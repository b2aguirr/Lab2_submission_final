-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     May 1 2019 17:43:45

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "latticehx1k" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of latticehx1k
entity latticehx1k is
port (
    led : out std_logic_vector(4 downto 0);
    to_ir : out std_logic;
    test2 : out std_logic;
    sd : out std_logic;
    test1 : out std_logic;
    o_serial_data : out std_logic;
    from_pc : in std_logic;
    test3 : out std_logic;
    clk_in : in std_logic);
end latticehx1k;

-- Architecture of latticehx1k
-- View name is \INTERFACE\
architecture \INTERFACE\ of latticehx1k is

signal \N__7037\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7026\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6983\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6974\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6938\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6929\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6908\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6905\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6867\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6823\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6795\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6793\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6787\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6763\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6749\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6739\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6711\ : std_logic;
signal \N__6708\ : std_logic;
signal \N__6705\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6663\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6603\ : std_logic;
signal \N__6600\ : std_logic;
signal \N__6597\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6534\ : std_logic;
signal \N__6531\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6510\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6474\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6438\ : std_logic;
signal \N__6431\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6413\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6360\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6354\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6340\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6333\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6309\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6291\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6186\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6072\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6041\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5996\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5917\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5812\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5785\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5716\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5409\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5382\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5198\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5140\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4768\ : std_logic;
signal \N__4765\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4417\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4294\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4285\ : std_logic;
signal \N__4282\ : std_logic;
signal \N__4279\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4230\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4219\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4186\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4181\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4123\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4120\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4114\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4089\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4074\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4060\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4030\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4027\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4015\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4003\ : std_logic;
signal \N__3994\ : std_logic;
signal \N__3991\ : std_logic;
signal \N__3988\ : std_logic;
signal \N__3987\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3985\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3975\ : std_logic;
signal \N__3970\ : std_logic;
signal \N__3969\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3967\ : std_logic;
signal \N__3964\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3949\ : std_logic;
signal \N__3946\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3941\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3937\ : std_logic;
signal \N__3934\ : std_logic;
signal \N__3929\ : std_logic;
signal \N__3928\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3922\ : std_logic;
signal \N__3919\ : std_logic;
signal \N__3916\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3908\ : std_logic;
signal \N__3907\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3905\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3899\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3856\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3853\ : std_logic;
signal \N__3852\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3850\ : std_logic;
signal \N__3849\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3844\ : std_logic;
signal \N__3841\ : std_logic;
signal \N__3838\ : std_logic;
signal \N__3835\ : std_logic;
signal \N__3832\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3802\ : std_logic;
signal \N__3799\ : std_logic;
signal \N__3796\ : std_logic;
signal \N__3793\ : std_logic;
signal \N__3790\ : std_logic;
signal \N__3787\ : std_logic;
signal \N__3784\ : std_logic;
signal \N__3781\ : std_logic;
signal \N__3778\ : std_logic;
signal \N__3775\ : std_logic;
signal \N__3772\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3766\ : std_logic;
signal \N__3763\ : std_logic;
signal \N__3760\ : std_logic;
signal \N__3757\ : std_logic;
signal \N__3754\ : std_logic;
signal \N__3751\ : std_logic;
signal \N__3748\ : std_logic;
signal \N__3745\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3733\ : std_logic;
signal \N__3730\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3726\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3718\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3706\ : std_logic;
signal \N__3705\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3703\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3690\ : std_logic;
signal \N__3687\ : std_logic;
signal \N__3684\ : std_logic;
signal \N__3679\ : std_logic;
signal \N__3676\ : std_logic;
signal \N__3673\ : std_logic;
signal \N__3672\ : std_logic;
signal \N__3669\ : std_logic;
signal \N__3668\ : std_logic;
signal \N__3665\ : std_logic;
signal \N__3662\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3653\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3647\ : std_logic;
signal \N__3642\ : std_logic;
signal \N__3637\ : std_logic;
signal \N__3634\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3627\ : std_logic;
signal \N__3624\ : std_logic;
signal \N__3621\ : std_logic;
signal \N__3616\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3607\ : std_logic;
signal \N__3604\ : std_logic;
signal \N__3601\ : std_logic;
signal \N__3598\ : std_logic;
signal \N__3595\ : std_logic;
signal \N__3592\ : std_logic;
signal \N__3589\ : std_logic;
signal \N__3586\ : std_logic;
signal \N__3583\ : std_logic;
signal \N__3580\ : std_logic;
signal \N__3579\ : std_logic;
signal \N__3576\ : std_logic;
signal \N__3573\ : std_logic;
signal \N__3572\ : std_logic;
signal \N__3567\ : std_logic;
signal \N__3564\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3558\ : std_logic;
signal \N__3557\ : std_logic;
signal \N__3552\ : std_logic;
signal \N__3549\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3543\ : std_logic;
signal \N__3538\ : std_logic;
signal \N__3535\ : std_logic;
signal \N__3534\ : std_logic;
signal \N__3533\ : std_logic;
signal \N__3528\ : std_logic;
signal \N__3527\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3523\ : std_logic;
signal \N__3522\ : std_logic;
signal \N__3519\ : std_logic;
signal \N__3516\ : std_logic;
signal \N__3513\ : std_logic;
signal \N__3508\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3496\ : std_logic;
signal \N__3493\ : std_logic;
signal \N__3490\ : std_logic;
signal \N__3487\ : std_logic;
signal \N__3484\ : std_logic;
signal \N__3481\ : std_logic;
signal \N__3478\ : std_logic;
signal \N__3475\ : std_logic;
signal \N__3472\ : std_logic;
signal \N__3469\ : std_logic;
signal \N__3466\ : std_logic;
signal \N__3463\ : std_logic;
signal \N__3462\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3456\ : std_logic;
signal \N__3451\ : std_logic;
signal \N__3448\ : std_logic;
signal \N__3447\ : std_logic;
signal \N__3446\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3444\ : std_logic;
signal \N__3443\ : std_logic;
signal \N__3440\ : std_logic;
signal \N__3437\ : std_logic;
signal \N__3434\ : std_logic;
signal \N__3427\ : std_logic;
signal \N__3424\ : std_logic;
signal \N__3421\ : std_logic;
signal \N__3412\ : std_logic;
signal \N__3409\ : std_logic;
signal \N__3408\ : std_logic;
signal \N__3407\ : std_logic;
signal \N__3404\ : std_logic;
signal \N__3401\ : std_logic;
signal \N__3398\ : std_logic;
signal \N__3391\ : std_logic;
signal \N__3390\ : std_logic;
signal \N__3387\ : std_logic;
signal \N__3384\ : std_logic;
signal \N__3381\ : std_logic;
signal \N__3376\ : std_logic;
signal \N__3375\ : std_logic;
signal \N__3374\ : std_logic;
signal \N__3373\ : std_logic;
signal \N__3370\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3362\ : std_logic;
signal \N__3359\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3349\ : std_logic;
signal \N__3346\ : std_logic;
signal \N__3343\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3337\ : std_logic;
signal \N__3334\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3328\ : std_logic;
signal \N__3325\ : std_logic;
signal \N__3322\ : std_logic;
signal \N__3321\ : std_logic;
signal \N__3320\ : std_logic;
signal \N__3319\ : std_logic;
signal \N__3318\ : std_logic;
signal \N__3317\ : std_logic;
signal \N__3312\ : std_logic;
signal \N__3307\ : std_logic;
signal \N__3304\ : std_logic;
signal \N__3301\ : std_logic;
signal \N__3292\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3288\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3284\ : std_logic;
signal \N__3283\ : std_logic;
signal \N__3280\ : std_logic;
signal \N__3277\ : std_logic;
signal \N__3274\ : std_logic;
signal \N__3271\ : std_logic;
signal \N__3268\ : std_logic;
signal \N__3259\ : std_logic;
signal \N__3258\ : std_logic;
signal \N__3255\ : std_logic;
signal \N__3254\ : std_logic;
signal \N__3253\ : std_logic;
signal \N__3250\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3246\ : std_logic;
signal \N__3241\ : std_logic;
signal \N__3236\ : std_logic;
signal \N__3229\ : std_logic;
signal \N__3226\ : std_logic;
signal \N__3223\ : std_logic;
signal \N__3220\ : std_logic;
signal \N__3217\ : std_logic;
signal \N__3214\ : std_logic;
signal \N__3213\ : std_logic;
signal \N__3212\ : std_logic;
signal \N__3211\ : std_logic;
signal \N__3208\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3200\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3192\ : std_logic;
signal \N__3191\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3185\ : std_logic;
signal \N__3182\ : std_logic;
signal \N__3175\ : std_logic;
signal \N__3172\ : std_logic;
signal \N__3169\ : std_logic;
signal \N__3166\ : std_logic;
signal \N__3163\ : std_logic;
signal \N__3160\ : std_logic;
signal \N__3157\ : std_logic;
signal \N__3154\ : std_logic;
signal \N__3151\ : std_logic;
signal \N__3148\ : std_logic;
signal \N__3145\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3133\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3129\ : std_logic;
signal \N__3126\ : std_logic;
signal \N__3123\ : std_logic;
signal \N__3120\ : std_logic;
signal \N__3119\ : std_logic;
signal \N__3116\ : std_logic;
signal \N__3113\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3107\ : std_logic;
signal \N__3104\ : std_logic;
signal \N__3099\ : std_logic;
signal \N__3094\ : std_logic;
signal \N__3091\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3085\ : std_logic;
signal \N__3082\ : std_logic;
signal \N__3079\ : std_logic;
signal \N__3076\ : std_logic;
signal \N__3073\ : std_logic;
signal \N__3070\ : std_logic;
signal \N__3067\ : std_logic;
signal \N__3064\ : std_logic;
signal \N__3061\ : std_logic;
signal \N__3058\ : std_logic;
signal \N__3055\ : std_logic;
signal \N__3052\ : std_logic;
signal \N__3049\ : std_logic;
signal \N__3046\ : std_logic;
signal \N__3043\ : std_logic;
signal \N__3040\ : std_logic;
signal \N__3037\ : std_logic;
signal \N__3034\ : std_logic;
signal \N__3031\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3022\ : std_logic;
signal \N__3019\ : std_logic;
signal \N__3016\ : std_logic;
signal \N__3013\ : std_logic;
signal \N__3010\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3004\ : std_logic;
signal \N__3001\ : std_logic;
signal \N__2998\ : std_logic;
signal \N__2995\ : std_logic;
signal \N__2992\ : std_logic;
signal \N__2989\ : std_logic;
signal \N__2986\ : std_logic;
signal \N__2983\ : std_logic;
signal \N__2980\ : std_logic;
signal \N__2977\ : std_logic;
signal \N__2974\ : std_logic;
signal \N__2971\ : std_logic;
signal \N__2970\ : std_logic;
signal \N__2967\ : std_logic;
signal \N__2964\ : std_logic;
signal \N__2959\ : std_logic;
signal \N__2956\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2950\ : std_logic;
signal \N__2947\ : std_logic;
signal \N__2944\ : std_logic;
signal \N__2941\ : std_logic;
signal \N__2938\ : std_logic;
signal \N__2935\ : std_logic;
signal \N__2932\ : std_logic;
signal \N__2929\ : std_logic;
signal \N__2926\ : std_logic;
signal \N__2923\ : std_logic;
signal \N__2920\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2914\ : std_logic;
signal \N__2911\ : std_logic;
signal \N__2908\ : std_logic;
signal \N__2905\ : std_logic;
signal \N__2902\ : std_logic;
signal \N__2899\ : std_logic;
signal \N__2896\ : std_logic;
signal \N__2893\ : std_logic;
signal \N__2892\ : std_logic;
signal \N__2889\ : std_logic;
signal \N__2886\ : std_logic;
signal \N__2881\ : std_logic;
signal \N__2878\ : std_logic;
signal \N__2875\ : std_logic;
signal \N__2872\ : std_logic;
signal \N__2871\ : std_logic;
signal \N__2868\ : std_logic;
signal \N__2865\ : std_logic;
signal \N__2860\ : std_logic;
signal \N__2857\ : std_logic;
signal \N__2854\ : std_logic;
signal \N__2851\ : std_logic;
signal \N__2848\ : std_logic;
signal \N__2845\ : std_logic;
signal \N__2842\ : std_logic;
signal \N__2839\ : std_logic;
signal \N__2838\ : std_logic;
signal \N__2835\ : std_logic;
signal \N__2832\ : std_logic;
signal \N__2829\ : std_logic;
signal \N__2826\ : std_logic;
signal \N__2823\ : std_logic;
signal \N__2818\ : std_logic;
signal \N__2815\ : std_logic;
signal \N__2812\ : std_logic;
signal \N__2809\ : std_logic;
signal \N__2806\ : std_logic;
signal \N__2803\ : std_logic;
signal \N__2800\ : std_logic;
signal \N__2797\ : std_logic;
signal \N__2794\ : std_logic;
signal \N__2791\ : std_logic;
signal \N__2788\ : std_logic;
signal \N__2785\ : std_logic;
signal \N__2782\ : std_logic;
signal \N__2779\ : std_logic;
signal \N__2776\ : std_logic;
signal \N__2773\ : std_logic;
signal \N__2770\ : std_logic;
signal \N__2767\ : std_logic;
signal \N__2764\ : std_logic;
signal \N__2761\ : std_logic;
signal \N__2758\ : std_logic;
signal \N__2755\ : std_logic;
signal \N__2752\ : std_logic;
signal \N__2749\ : std_logic;
signal \N__2746\ : std_logic;
signal \VCCG0\ : std_logic;
signal clk_in_c : std_logic;
signal clk : std_logic;
signal \GNDG0\ : std_logic;
signal \uart_RXD\ : std_logic;
signal o_serial_data_c : std_logic;
signal \bfn_6_11_0_\ : std_logic;
signal \Glue_Lab2.reset_count_cry_0\ : std_logic;
signal \Glue_Lab2.reset_count_cry_1\ : std_logic;
signal \Glue_Lab2.reset_count_cry_2\ : std_logic;
signal \Glue_Lab2.reset_count_cry_3\ : std_logic;
signal \Glue_Lab2.reset_count_cry_1_THRU_CO\ : std_logic;
signal \Glue_Lab2.reset_countZ0Z_2\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_1\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_0\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_2\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_3\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_4\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_5\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_7\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_6\ : std_logic;
signal \Glue_Lab2.reset_count_cry_2_THRU_CO\ : std_logic;
signal \Glue_Lab2.reset_countZ0Z_3\ : std_logic;
signal \Glue_Lab2.reset_count_cry_0_THRU_CO\ : std_logic;
signal \Glue_Lab2.reset_countZ0Z_1\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counter_0_1_5_cascade_\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_ac0_7\ : std_logic;
signal \buart.Z_rx.ser_clk_2_cascade_\ : std_logic;
signal \Glue_Lab2.reset_countZ0Z_0\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_4\ : std_logic;
signal \Lab_UT.sDelay.delayRegZ0Z_0\ : std_logic;
signal \Gl_tx_data_0\ : std_logic;
signal \Lab_UT.S_m_bmZ0Z_3_cascade_\ : std_logic;
signal led_c_3 : std_logic;
signal \led_c_3_cascade_\ : std_logic;
signal \Gl_tx_data_3\ : std_logic;
signal \Lab_UT.S_m_bm_N_3LZ0Z3\ : std_logic;
signal \Lab_UT.g0_0_a3_0Z0Z_0_cascade_\ : std_logic;
signal \Lab_UT_C_out41_1_cascade_\ : std_logic;
signal \Gl_tx_data_5\ : std_logic;
signal \Lab_UT.N_6_0\ : std_logic;
signal \Lab_UT.g0_0_a3Z0Z_0_cascade_\ : std_logic;
signal \Lab_UT.g0_1Z0Z_0\ : std_logic;
signal \Lab_UT.N_6\ : std_logic;
signal \Lab_UT.S_0_s_axbZ0Z3_cascade_\ : std_logic;
signal \Lab_UT.S_m_amZ0Z_3\ : std_logic;
signal \Lab_UT.g1_0_0\ : std_logic;
signal \Lab_UT.S_m_bm_N_6LZ0Z10\ : std_logic;
signal \Glue_Lab2.g0_9_0_cascade_\ : std_logic;
signal \Glue_Lab2.reset_counte_0_1\ : std_logic;
signal \Glue_Lab2.g0_7_0\ : std_logic;
signal \buart.Z_rx.bitcountlde_0_cascade_\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \buart.Z_rx.N_29_0_i_cascade_\ : std_logic;
signal \buart.Z_rx.bitcount_lm_0\ : std_logic;
signal \Glue_Lab2.de0.g0_5_0\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_0\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_1\ : std_logic;
signal \Glue_Lab2.de0.g0_5_2_cascade_\ : std_logic;
signal \Glue_Lab2.g0_9_2_cascade_\ : std_logic;
signal \Glue_Lab2.g0_7_2\ : std_logic;
signal \Glue_Lab2.reset_counte_0_3\ : std_logic;
signal \buart.Z_rx.bitcount_RNIMK771_0Z0Z_4_cascade_\ : std_logic;
signal \bu_rx_data_rdy_cascade_\ : std_logic;
signal \Glue_Lab2.i_rst_char_detected\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_4\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_5\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_3\ : std_logic;
signal \buart.Z_rx.un1_sample_0\ : std_logic;
signal \buart.Z_rx.ser_clk_2_0_cascade_\ : std_logic;
signal \Glue_Lab2.de0.un2_de_hexplus_3_xZ0Z0_cascade_\ : std_logic;
signal \Glue_Lab2.de0.un2_de_hexplus_3_cascade_\ : std_logic;
signal \Glue_Lab2.is_hexplus_cascade_\ : std_logic;
signal \Gl_tx_data_4\ : std_logic;
signal \buart.Z_rx.ser_clk_2\ : std_logic;
signal \buart.Z_rx.ser_clk_2_0\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_2\ : std_logic;
signal \Glue_Lab2.gl_fsm.N_14_cascade_\ : std_logic;
signal \Glue_Lab2_gl_fsm_state_0\ : std_logic;
signal \Lab_UT.C_out41_0\ : std_logic;
signal \led_c_0_4_cascade_\ : std_logic;
signal \Gl_tx_data_6\ : std_logic;
signal \Lab_UT.S_m_bm_N_2LZ0Z1\ : std_logic;
signal led_c_0 : std_logic;
signal \Lab_UT.S_1_ac0_1_0Z0Z_0\ : std_logic;
signal \Lab_UT.S_1_axbZ0Z1_cascade_\ : std_logic;
signal \Lab_UT.g1Z0Z_0\ : std_logic;
signal \Lab_UT.S_0_s_c2_0_cascade_\ : std_logic;
signal \Lab_UT.S_0_s_ac0_5_0_1\ : std_logic;
signal \Lab_UT.gZ0Z1\ : std_logic;
signal \Glue_Lab2_Gl_r2_fast_0\ : std_logic;
signal \Glue_Lab2_Gl_r1_fast_0\ : std_logic;
signal \Lab_UT.S_m_bm_N_5LZ0Z7\ : std_logic;
signal \Gl_r1_2_rep1\ : std_logic;
signal \Gl_r2_2_rep1\ : std_logic;
signal \Lab_UT.g0_4Z0Z_0\ : std_logic;
signal \Glue_Lab2.Gl_r17_0_i\ : std_logic;
signal \Lab_UT.g0_1_0_0\ : std_logic;
signal \Glue_Lab2.Gl_r27_0_i\ : std_logic;
signal \Lab_UT.g0_4_0_0\ : std_logic;
signal \Lab_UT.S_0_s_c2_1_cascade_\ : std_logic;
signal \Lab_UT.S_0_s_ac0_5_0_2\ : std_logic;
signal \Lab_UT_g1_1\ : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal \buart.Z_rx.bitcount_cry_0\ : std_logic;
signal \buart.Z_rx.bitcount_cry_1\ : std_logic;
signal \buart.Z_rx.bitcount_cry_2\ : std_logic;
signal \buart.Z_rx.bitcount_cry_3\ : std_logic;
signal \buart.Z_rx.bitcount_lm_4\ : std_logic;
signal \buart.Z_rx.bitcount_cry_0_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcount_cry_2_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcount_lm_3_cascade_\ : std_logic;
signal \buart__rx_bitcount_4\ : std_logic;
signal \buart__rx_bitcount_3\ : std_logic;
signal \buart.Z_rx.bitcount_RNIMK771Z0Z_4_cascade_\ : std_logic;
signal \buart.Z_rx.idle\ : std_logic;
signal \buart.Z_rx.idle_cascade_\ : std_logic;
signal \buart.Z_rx.hhZ0Z_0\ : std_logic;
signal \buart.Z_rx.startbit_cascade_\ : std_logic;
signal \buart.Z_rx.bitcount_lm_1\ : std_logic;
signal \buart__rx_bitcount_1\ : std_logic;
signal \buart.Z_rx.bitcount_cry_1_THRU_CO\ : std_logic;
signal \buart.Z_rx.N_29_0_i\ : std_logic;
signal \buart.Z_rx.bitcountlde_0\ : std_logic;
signal \buart.Z_rx.bitcount_lm_2_cascade_\ : std_logic;
signal \buart.Z_rx.startbit\ : std_logic;
signal \buart__rx_bitcount_2\ : std_logic;
signal \Glue_Lab2.g0_8_2\ : std_logic;
signal \Glue_Lab2.de0.un2_de_hexplusZ0Z_2\ : std_logic;
signal \Glue_Lab2.de0.un1_charDataZ0\ : std_logic;
signal \buart__rx_shifter_fast_5\ : std_logic;
signal \buart.Z_rx.hhZ0Z_1\ : std_logic;
signal \Glue_Lab2.g0_8_0\ : std_logic;
signal \Glue_Lab2.de0.de_escZ0Z_3\ : std_logic;
signal \Glue_Lab2.gl_fsm.enOp_0_a2_1\ : std_logic;
signal \Glue_Lab2.gl_fsm.enOp_0_a2Z0Z_4\ : std_logic;
signal bu_rx_data_rdy : std_logic;
signal \Glue_Lab2.Gl_r1_2_1_cascade_\ : std_logic;
signal \Glue_Lab2.Gl_r1_2_2_cascade_\ : std_logic;
signal \Lab_UT.g0Z0Z_1\ : std_logic;
signal \Glue_Lab2.enOp\ : std_logic;
signal \Gl_tx_data_2\ : std_logic;
signal \Glue_Lab2_gl_fsm_state_1\ : std_logic;
signal \Glue_Lab2.gl_fsm.enOp_0_a2_2\ : std_logic;
signal \Glue_Lab2.Gl_subtract_1_cascade_\ : std_logic;
signal \Lab_UT.S_0_s_axbZ0Z3\ : std_logic;
signal \Lab_UT.S_0_s_cZ0Z2\ : std_logic;
signal \Lab_UT.S_m_amZ0Z_2_cascade_\ : std_logic;
signal led_c_2 : std_logic;
signal \Gl_r1_0\ : std_logic;
signal \Gl_r2_1\ : std_logic;
signal \Gl_r2_0\ : std_logic;
signal \Gl_r1_1\ : std_logic;
signal \Lab_UT.S_m_amZ0Z_1\ : std_logic;
signal \Lab_UT.S_m_bmZ0Z_1_cascade_\ : std_logic;
signal led_c_1 : std_logic;
signal \led_c_1_cascade_\ : std_logic;
signal \Gl_tx_data_1\ : std_logic;
signal \Gl_r2_fast_2\ : std_logic;
signal \Gl_r1_fast_2\ : std_logic;
signal \Lab_UT.S_m_bm_1Z0Z_2\ : std_logic;
signal \Lab_UT.S_m_bmZ0Z_2\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_c5_cascade_\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_c5\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_5\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_6\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_1\ : std_logic;
signal \buart.Z_tx.Z_baudgen.ser_clk_sx_cascade_\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_0\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counter_RNIES38_0Z0Z_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un1_bitcount_c2_1\ : std_logic;
signal \buart.Z_tx.bitcount_RNIBADLZ0Z_1_cascade_\ : std_logic;
signal \buart.Z_tx.counter_RNIVE1P1_4_cascade_\ : std_logic;
signal \buart.Z_tx.un1_bitcount_c2\ : std_logic;
signal \buart.Z_tx.uart_busy_0_0\ : std_logic;
signal \buart.Z_tx.uart_busy_0_0_cascade_\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_2\ : std_logic;
signal \buart.Z_tx.un1_bitcount_c3_cascade_\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_3\ : std_logic;
signal \buart.Z_tx.un1_uart_wr_i_0_i_sx\ : std_logic;
signal \Glue_Lab2.is_hexplus\ : std_logic;
signal \buart.Z_tx.un1_bitcount_c1_cascade_\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_1\ : std_logic;
signal \buart.Z_tx.counter_RNIVE1P1_4\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_0\ : std_logic;
signal \Glue_Lab2.de0.de_escZ0Z_4\ : std_logic;
signal \Glue_Lab2.de0.g0_5_1_cascade_\ : std_logic;
signal \Glue_Lab2.g0_9_1_cascade_\ : std_logic;
signal \Glue_Lab2.g0_7_1\ : std_logic;
signal \Glue_Lab2.reset_counte_0_2\ : std_logic;
signal bu_rx_data_4 : std_logic;
signal \buart__rx_bitcount_0\ : std_logic;
signal \Glue_Lab2.de0.g0Z0Z_5_cascade_\ : std_logic;
signal bu_rx_data_0 : std_logic;
signal \Glue_Lab2.reset_countZ0Z_4\ : std_logic;
signal \Glue_Lab2.g0_9_cascade_\ : std_logic;
signal \Glue_Lab2.g0_7\ : std_logic;
signal \Glue_Lab2.reset_counte_0_0\ : std_logic;
signal bu_rx_data_2 : std_logic;
signal bu_rx_data_6 : std_logic;
signal \buart__rx_shifter_fast_4\ : std_logic;
signal \buart.Z_rx.sample\ : std_logic;
signal \Glue_Lab2_Gl_Op_0\ : std_logic;
signal \Glue_Lab2_Gl_Op_3\ : std_logic;
signal \Glue_Lab2_Gl_Op_1\ : std_logic;
signal \Glue_Lab2_Gl_Op_5\ : std_logic;
signal \Glue_Lab2.g0_0_1_0_cascade_\ : std_logic;
signal \Glue_Lab2_Gl_Op_2\ : std_logic;
signal \Glue_Lab2.Gl_subtract_0\ : std_logic;
signal \Gl_r1_2\ : std_logic;
signal \Gl_r2_2\ : std_logic;
signal \Gl_r1_3\ : std_logic;
signal \Lab_UT.S_1_c3_d\ : std_logic;
signal \Lab_UT.S_1_c3_cZ0_cascade_\ : std_logic;
signal \Gl_r2_3\ : std_logic;
signal \Lab_UT.S_0_s_ac0_5_0Z0Z_0\ : std_logic;
signal \Lab_UT.S_0_s_ac0_5_dZ0\ : std_logic;
signal \Lab_UT.C_out41_cascade_\ : std_logic;
signal \Gl_subtract\ : std_logic;
signal led_c_4 : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_2\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_c2\ : std_logic;
signal \buart.Z_tx.ser_clk\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_3\ : std_logic;
signal \Gl_tx_data_rdy\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_8\ : std_logic;
signal \buart.Z_tx.un1_uart_wr_i_0_i\ : std_logic;
signal \Glue_Lab2.g0_8\ : std_logic;
signal bu_rx_data_7 : std_logic;
signal bu_rx_data_3 : std_logic;
signal bu_rx_data_5 : std_logic;
signal bu_rx_data_1 : std_logic;
signal \Glue_Lab2.g0_8_1\ : std_logic;
signal \Lab_UT.sDelay.delayRegZ0Z_1\ : std_logic;
signal \Lab_UT.sDelay.delayRegZ0Z_2\ : std_logic;
signal \Lab_UT.sDelay.delayRegZ0Z_3\ : std_logic;
signal \Gl_rst\ : std_logic;
signal \L2_adder_rdy\ : std_logic;
signal clk_g : std_logic;
signal \_gnd_net_\ : std_logic;

signal led_wire : std_logic_vector(4 downto 0);
signal test1_wire : std_logic;
signal from_pc_wire : std_logic;
signal sd_wire : std_logic;
signal clk_in_wire : std_logic;
signal test3_wire : std_logic;
signal to_ir_wire : std_logic;
signal o_serial_data_wire : std_logic;
signal test2_wire : std_logic;
signal \ice_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    led <= led_wire;
    test1 <= test1_wire;
    from_pc_wire <= from_pc;
    sd <= sd_wire;
    clk_in_wire <= clk_in;
    test3 <= test3_wire;
    to_ir <= to_ir_wire;
    o_serial_data <= o_serial_data_wire;
    test2 <= test2_wire;
    \ice_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \ice_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "100",
            DIVF => "0111111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => clk,
            REFERENCECLK => \N__2806\,
            RESETB => \N__3133\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \ice_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \led_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7037\,
            DIN => \N__7036\,
            DOUT => \N__7035\,
            PACKAGEPIN => led_wire(0)
        );

    \led_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7037\,
            PADOUT => \N__7036\,
            PADIN => \N__7035\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3469\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \test1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7028\,
            DIN => \N__7027\,
            DOUT => \N__7026\,
            PACKAGEPIN => test1_wire
        );

    \test1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7028\,
            PADOUT => \N__7027\,
            PADIN => \N__7026\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Z_rcxd.Z_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7019\,
            DIN => \N__7018\,
            DOUT => \N__7017\,
            PACKAGEPIN => from_pc_wire
        );

    \Z_rcxd.Z_io_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__7019\,
            PADOUT => \N__7018\,
            PADIN => \N__7017\,
            CLOCKENABLE => 'H',
            DOUT1 => \GNDG0\,
            OUTPUTENABLE => '0',
            DIN0 => \uart_RXD\,
            DOUT0 => \GNDG0\,
            INPUTCLK => \N__6162\,
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \sd_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7010\,
            DIN => \N__7009\,
            DOUT => \N__7008\,
            PACKAGEPIN => sd_wire
        );

    \sd_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7010\,
            PADOUT => \N__7009\,
            PADIN => \N__7008\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clk_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7001\,
            DIN => \N__7000\,
            DOUT => \N__6999\,
            PACKAGEPIN => clk_in_wire
        );

    \clk_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7001\,
            PADOUT => \N__7000\,
            PADIN => \N__6999\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => clk_in_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6992\,
            DIN => \N__6991\,
            DOUT => \N__6990\,
            PACKAGEPIN => led_wire(2)
        );

    \led_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6992\,
            PADOUT => \N__6991\,
            PADIN => \N__6990\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4621\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6983\,
            DIN => \N__6982\,
            DOUT => \N__6981\,
            PACKAGEPIN => led_wire(4)
        );

    \led_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6983\,
            PADOUT => \N__6982\,
            PADIN => \N__6981\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5542\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \test3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6974\,
            DIN => \N__6973\,
            DOUT => \N__6972\,
            PACKAGEPIN => test3_wire
        );

    \test3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6974\,
            PADOUT => \N__6973\,
            PADIN => \N__6972\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \to_ir_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6965\,
            DIN => \N__6964\,
            DOUT => \N__6963\,
            PACKAGEPIN => to_ir_wire
        );

    \to_ir_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6965\,
            PADOUT => \N__6964\,
            PADIN => \N__6963\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6956\,
            DIN => \N__6955\,
            DOUT => \N__6954\,
            PACKAGEPIN => led_wire(1)
        );

    \led_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6956\,
            PADOUT => \N__6955\,
            PADIN => \N__6954\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4342\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6947\,
            DIN => \N__6946\,
            DOUT => \N__6945\,
            PACKAGEPIN => led_wire(3)
        );

    \led_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6947\,
            PADOUT => \N__6946\,
            PADIN => \N__6945\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3034\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_serial_data_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6938\,
            DIN => \N__6937\,
            DOUT => \N__6936\,
            PACKAGEPIN => o_serial_data_wire
        );

    \o_serial_data_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6938\,
            PADOUT => \N__6937\,
            PADIN => \N__6936\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2761\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \test2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6929\,
            DIN => \N__6928\,
            DOUT => \N__6927\,
            PACKAGEPIN => test2_wire
        );

    \test2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6929\,
            PADOUT => \N__6928\,
            PADIN => \N__6927\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1620\ : InMux
    port map (
            O => \N__6910\,
            I => \N__6900\
        );

    \I__1619\ : InMux
    port map (
            O => \N__6909\,
            I => \N__6900\
        );

    \I__1618\ : InMux
    port map (
            O => \N__6908\,
            I => \N__6891\
        );

    \I__1617\ : InMux
    port map (
            O => \N__6907\,
            I => \N__6891\
        );

    \I__1616\ : InMux
    port map (
            O => \N__6906\,
            I => \N__6891\
        );

    \I__1615\ : InMux
    port map (
            O => \N__6905\,
            I => \N__6891\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__6900\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_2\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__6891\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_2\
        );

    \I__1612\ : CascadeMux
    port map (
            O => \N__6886\,
            I => \N__6882\
        );

    \I__1611\ : CascadeMux
    port map (
            O => \N__6885\,
            I => \N__6878\
        );

    \I__1610\ : InMux
    port map (
            O => \N__6882\,
            I => \N__6872\
        );

    \I__1609\ : InMux
    port map (
            O => \N__6881\,
            I => \N__6872\
        );

    \I__1608\ : InMux
    port map (
            O => \N__6878\,
            I => \N__6867\
        );

    \I__1607\ : InMux
    port map (
            O => \N__6877\,
            I => \N__6867\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__6872\,
            I => \N__6864\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__6867\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_c2\
        );

    \I__1604\ : Odrv4
    port map (
            O => \N__6864\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_c2\
        );

    \I__1603\ : InMux
    port map (
            O => \N__6859\,
            I => \N__6850\
        );

    \I__1602\ : InMux
    port map (
            O => \N__6858\,
            I => \N__6850\
        );

    \I__1601\ : InMux
    port map (
            O => \N__6857\,
            I => \N__6845\
        );

    \I__1600\ : InMux
    port map (
            O => \N__6856\,
            I => \N__6840\
        );

    \I__1599\ : InMux
    port map (
            O => \N__6855\,
            I => \N__6840\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__6850\,
            I => \N__6837\
        );

    \I__1597\ : InMux
    port map (
            O => \N__6849\,
            I => \N__6832\
        );

    \I__1596\ : InMux
    port map (
            O => \N__6848\,
            I => \N__6832\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__6845\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__6840\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__1593\ : Odrv4
    port map (
            O => \N__6837\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__6832\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__1591\ : CascadeMux
    port map (
            O => \N__6823\,
            I => \N__6817\
        );

    \I__1590\ : CascadeMux
    port map (
            O => \N__6822\,
            I => \N__6814\
        );

    \I__1589\ : InMux
    port map (
            O => \N__6821\,
            I => \N__6810\
        );

    \I__1588\ : InMux
    port map (
            O => \N__6820\,
            I => \N__6801\
        );

    \I__1587\ : InMux
    port map (
            O => \N__6817\,
            I => \N__6801\
        );

    \I__1586\ : InMux
    port map (
            O => \N__6814\,
            I => \N__6801\
        );

    \I__1585\ : InMux
    port map (
            O => \N__6813\,
            I => \N__6801\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__6810\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_3\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__6801\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_3\
        );

    \I__1582\ : InMux
    port map (
            O => \N__6796\,
            I => \N__6782\
        );

    \I__1581\ : InMux
    port map (
            O => \N__6795\,
            I => \N__6765\
        );

    \I__1580\ : InMux
    port map (
            O => \N__6794\,
            I => \N__6765\
        );

    \I__1579\ : InMux
    port map (
            O => \N__6793\,
            I => \N__6765\
        );

    \I__1578\ : InMux
    port map (
            O => \N__6792\,
            I => \N__6765\
        );

    \I__1577\ : InMux
    port map (
            O => \N__6791\,
            I => \N__6765\
        );

    \I__1576\ : InMux
    port map (
            O => \N__6790\,
            I => \N__6765\
        );

    \I__1575\ : InMux
    port map (
            O => \N__6789\,
            I => \N__6765\
        );

    \I__1574\ : InMux
    port map (
            O => \N__6788\,
            I => \N__6765\
        );

    \I__1573\ : InMux
    port map (
            O => \N__6787\,
            I => \N__6754\
        );

    \I__1572\ : InMux
    port map (
            O => \N__6786\,
            I => \N__6754\
        );

    \I__1571\ : InMux
    port map (
            O => \N__6785\,
            I => \N__6754\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__6782\,
            I => \N__6749\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__6765\,
            I => \N__6749\
        );

    \I__1568\ : InMux
    port map (
            O => \N__6764\,
            I => \N__6746\
        );

    \I__1567\ : InMux
    port map (
            O => \N__6763\,
            I => \N__6739\
        );

    \I__1566\ : InMux
    port map (
            O => \N__6762\,
            I => \N__6739\
        );

    \I__1565\ : InMux
    port map (
            O => \N__6761\,
            I => \N__6739\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__6754\,
            I => \N__6736\
        );

    \I__1563\ : Odrv12
    port map (
            O => \N__6749\,
            I => \Gl_tx_data_rdy\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__6746\,
            I => \Gl_tx_data_rdy\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__6739\,
            I => \Gl_tx_data_rdy\
        );

    \I__1560\ : Odrv4
    port map (
            O => \N__6736\,
            I => \Gl_tx_data_rdy\
        );

    \I__1559\ : InMux
    port map (
            O => \N__6727\,
            I => \N__6724\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__6724\,
            I => \N__6721\
        );

    \I__1557\ : Span4Mux_h
    port map (
            O => \N__6721\,
            I => \N__6718\
        );

    \I__1556\ : Odrv4
    port map (
            O => \N__6718\,
            I => \buart.Z_tx.shifterZ0Z_8\
        );

    \I__1555\ : CEMux
    port map (
            O => \N__6715\,
            I => \N__6712\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__6712\,
            I => \N__6708\
        );

    \I__1553\ : CEMux
    port map (
            O => \N__6711\,
            I => \N__6705\
        );

    \I__1552\ : Span4Mux_h
    port map (
            O => \N__6708\,
            I => \N__6702\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__6705\,
            I => \N__6698\
        );

    \I__1550\ : Span4Mux_s1_h
    port map (
            O => \N__6702\,
            I => \N__6695\
        );

    \I__1549\ : CEMux
    port map (
            O => \N__6701\,
            I => \N__6692\
        );

    \I__1548\ : Odrv12
    port map (
            O => \N__6698\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i\
        );

    \I__1547\ : Odrv4
    port map (
            O => \N__6695\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__6692\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i\
        );

    \I__1545\ : InMux
    port map (
            O => \N__6685\,
            I => \N__6682\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__6682\,
            I => \Glue_Lab2.g0_8\
        );

    \I__1543\ : InMux
    port map (
            O => \N__6679\,
            I => \N__6676\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__6676\,
            I => \N__6669\
        );

    \I__1541\ : InMux
    port map (
            O => \N__6675\,
            I => \N__6666\
        );

    \I__1540\ : InMux
    port map (
            O => \N__6674\,
            I => \N__6663\
        );

    \I__1539\ : CascadeMux
    port map (
            O => \N__6673\,
            I => \N__6656\
        );

    \I__1538\ : CascadeMux
    port map (
            O => \N__6672\,
            I => \N__6653\
        );

    \I__1537\ : Span4Mux_s2_h
    port map (
            O => \N__6669\,
            I => \N__6650\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__6666\,
            I => \N__6647\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__6663\,
            I => \N__6644\
        );

    \I__1534\ : InMux
    port map (
            O => \N__6662\,
            I => \N__6639\
        );

    \I__1533\ : InMux
    port map (
            O => \N__6661\,
            I => \N__6639\
        );

    \I__1532\ : InMux
    port map (
            O => \N__6660\,
            I => \N__6630\
        );

    \I__1531\ : InMux
    port map (
            O => \N__6659\,
            I => \N__6630\
        );

    \I__1530\ : InMux
    port map (
            O => \N__6656\,
            I => \N__6630\
        );

    \I__1529\ : InMux
    port map (
            O => \N__6653\,
            I => \N__6630\
        );

    \I__1528\ : Odrv4
    port map (
            O => \N__6650\,
            I => bu_rx_data_7
        );

    \I__1527\ : Odrv12
    port map (
            O => \N__6647\,
            I => bu_rx_data_7
        );

    \I__1526\ : Odrv4
    port map (
            O => \N__6644\,
            I => bu_rx_data_7
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__6639\,
            I => bu_rx_data_7
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__6630\,
            I => bu_rx_data_7
        );

    \I__1523\ : InMux
    port map (
            O => \N__6619\,
            I => \N__6616\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__6616\,
            I => \N__6609\
        );

    \I__1521\ : InMux
    port map (
            O => \N__6615\,
            I => \N__6606\
        );

    \I__1520\ : InMux
    port map (
            O => \N__6614\,
            I => \N__6603\
        );

    \I__1519\ : InMux
    port map (
            O => \N__6613\,
            I => \N__6600\
        );

    \I__1518\ : InMux
    port map (
            O => \N__6612\,
            I => \N__6597\
        );

    \I__1517\ : Span4Mux_s1_v
    port map (
            O => \N__6609\,
            I => \N__6590\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__6606\,
            I => \N__6590\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__6603\,
            I => \N__6587\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__6600\,
            I => \N__6582\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__6597\,
            I => \N__6582\
        );

    \I__1512\ : InMux
    port map (
            O => \N__6596\,
            I => \N__6579\
        );

    \I__1511\ : CascadeMux
    port map (
            O => \N__6595\,
            I => \N__6573\
        );

    \I__1510\ : Span4Mux_v
    port map (
            O => \N__6590\,
            I => \N__6569\
        );

    \I__1509\ : Span4Mux_h
    port map (
            O => \N__6587\,
            I => \N__6566\
        );

    \I__1508\ : Span4Mux_s2_h
    port map (
            O => \N__6582\,
            I => \N__6563\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__6579\,
            I => \N__6560\
        );

    \I__1506\ : InMux
    port map (
            O => \N__6578\,
            I => \N__6555\
        );

    \I__1505\ : InMux
    port map (
            O => \N__6577\,
            I => \N__6555\
        );

    \I__1504\ : InMux
    port map (
            O => \N__6576\,
            I => \N__6548\
        );

    \I__1503\ : InMux
    port map (
            O => \N__6573\,
            I => \N__6548\
        );

    \I__1502\ : InMux
    port map (
            O => \N__6572\,
            I => \N__6548\
        );

    \I__1501\ : Odrv4
    port map (
            O => \N__6569\,
            I => bu_rx_data_3
        );

    \I__1500\ : Odrv4
    port map (
            O => \N__6566\,
            I => bu_rx_data_3
        );

    \I__1499\ : Odrv4
    port map (
            O => \N__6563\,
            I => bu_rx_data_3
        );

    \I__1498\ : Odrv4
    port map (
            O => \N__6560\,
            I => bu_rx_data_3
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__6555\,
            I => bu_rx_data_3
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__6548\,
            I => bu_rx_data_3
        );

    \I__1495\ : CascadeMux
    port map (
            O => \N__6535\,
            I => \N__6531\
        );

    \I__1494\ : CascadeMux
    port map (
            O => \N__6534\,
            I => \N__6525\
        );

    \I__1493\ : InMux
    port map (
            O => \N__6531\,
            I => \N__6520\
        );

    \I__1492\ : InMux
    port map (
            O => \N__6530\,
            I => \N__6520\
        );

    \I__1491\ : CascadeMux
    port map (
            O => \N__6529\,
            I => \N__6516\
        );

    \I__1490\ : CascadeMux
    port map (
            O => \N__6528\,
            I => \N__6513\
        );

    \I__1489\ : InMux
    port map (
            O => \N__6525\,
            I => \N__6510\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__6520\,
            I => \N__6507\
        );

    \I__1487\ : InMux
    port map (
            O => \N__6519\,
            I => \N__6502\
        );

    \I__1486\ : InMux
    port map (
            O => \N__6516\,
            I => \N__6499\
        );

    \I__1485\ : InMux
    port map (
            O => \N__6513\,
            I => \N__6496\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__6510\,
            I => \N__6491\
        );

    \I__1483\ : Span4Mux_v
    port map (
            O => \N__6507\,
            I => \N__6491\
        );

    \I__1482\ : InMux
    port map (
            O => \N__6506\,
            I => \N__6486\
        );

    \I__1481\ : InMux
    port map (
            O => \N__6505\,
            I => \N__6486\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__6502\,
            I => bu_rx_data_5
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__6499\,
            I => bu_rx_data_5
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__6496\,
            I => bu_rx_data_5
        );

    \I__1477\ : Odrv4
    port map (
            O => \N__6491\,
            I => bu_rx_data_5
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__6486\,
            I => bu_rx_data_5
        );

    \I__1475\ : InMux
    port map (
            O => \N__6475\,
            I => \N__6466\
        );

    \I__1474\ : InMux
    port map (
            O => \N__6474\,
            I => \N__6463\
        );

    \I__1473\ : InMux
    port map (
            O => \N__6473\,
            I => \N__6457\
        );

    \I__1472\ : InMux
    port map (
            O => \N__6472\,
            I => \N__6454\
        );

    \I__1471\ : CascadeMux
    port map (
            O => \N__6471\,
            I => \N__6451\
        );

    \I__1470\ : InMux
    port map (
            O => \N__6470\,
            I => \N__6447\
        );

    \I__1469\ : CascadeMux
    port map (
            O => \N__6469\,
            I => \N__6443\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__6466\,
            I => \N__6438\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__6463\,
            I => \N__6438\
        );

    \I__1466\ : InMux
    port map (
            O => \N__6462\,
            I => \N__6431\
        );

    \I__1465\ : InMux
    port map (
            O => \N__6461\,
            I => \N__6431\
        );

    \I__1464\ : InMux
    port map (
            O => \N__6460\,
            I => \N__6431\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__6457\,
            I => \N__6428\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__6454\,
            I => \N__6425\
        );

    \I__1461\ : InMux
    port map (
            O => \N__6451\,
            I => \N__6422\
        );

    \I__1460\ : InMux
    port map (
            O => \N__6450\,
            I => \N__6419\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__6447\,
            I => \N__6416\
        );

    \I__1458\ : InMux
    port map (
            O => \N__6446\,
            I => \N__6413\
        );

    \I__1457\ : InMux
    port map (
            O => \N__6443\,
            I => \N__6410\
        );

    \I__1456\ : Span4Mux_v
    port map (
            O => \N__6438\,
            I => \N__6399\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__6431\,
            I => \N__6399\
        );

    \I__1454\ : Span4Mux_s0_h
    port map (
            O => \N__6428\,
            I => \N__6399\
        );

    \I__1453\ : Span4Mux_v
    port map (
            O => \N__6425\,
            I => \N__6399\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__6422\,
            I => \N__6399\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__6419\,
            I => bu_rx_data_1
        );

    \I__1450\ : Odrv12
    port map (
            O => \N__6416\,
            I => bu_rx_data_1
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__6413\,
            I => bu_rx_data_1
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__6410\,
            I => bu_rx_data_1
        );

    \I__1447\ : Odrv4
    port map (
            O => \N__6399\,
            I => bu_rx_data_1
        );

    \I__1446\ : InMux
    port map (
            O => \N__6388\,
            I => \N__6385\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__6385\,
            I => \Glue_Lab2.g0_8_1\
        );

    \I__1444\ : InMux
    port map (
            O => \N__6382\,
            I => \N__6379\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__6379\,
            I => \N__6376\
        );

    \I__1442\ : Odrv12
    port map (
            O => \N__6376\,
            I => \Lab_UT.sDelay.delayRegZ0Z_1\
        );

    \I__1441\ : InMux
    port map (
            O => \N__6373\,
            I => \N__6370\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__6370\,
            I => \Lab_UT.sDelay.delayRegZ0Z_2\
        );

    \I__1439\ : InMux
    port map (
            O => \N__6367\,
            I => \N__6364\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__6364\,
            I => \Lab_UT.sDelay.delayRegZ0Z_3\
        );

    \I__1437\ : CascadeMux
    port map (
            O => \N__6361\,
            I => \N__6349\
        );

    \I__1436\ : CascadeMux
    port map (
            O => \N__6360\,
            I => \N__6345\
        );

    \I__1435\ : CascadeMux
    port map (
            O => \N__6359\,
            I => \N__6340\
        );

    \I__1434\ : InMux
    port map (
            O => \N__6358\,
            I => \N__6333\
        );

    \I__1433\ : InMux
    port map (
            O => \N__6357\,
            I => \N__6324\
        );

    \I__1432\ : InMux
    port map (
            O => \N__6356\,
            I => \N__6324\
        );

    \I__1431\ : InMux
    port map (
            O => \N__6355\,
            I => \N__6324\
        );

    \I__1430\ : InMux
    port map (
            O => \N__6354\,
            I => \N__6324\
        );

    \I__1429\ : InMux
    port map (
            O => \N__6353\,
            I => \N__6319\
        );

    \I__1428\ : InMux
    port map (
            O => \N__6352\,
            I => \N__6319\
        );

    \I__1427\ : InMux
    port map (
            O => \N__6349\,
            I => \N__6314\
        );

    \I__1426\ : InMux
    port map (
            O => \N__6348\,
            I => \N__6314\
        );

    \I__1425\ : InMux
    port map (
            O => \N__6345\,
            I => \N__6301\
        );

    \I__1424\ : InMux
    port map (
            O => \N__6344\,
            I => \N__6301\
        );

    \I__1423\ : InMux
    port map (
            O => \N__6343\,
            I => \N__6292\
        );

    \I__1422\ : InMux
    port map (
            O => \N__6340\,
            I => \N__6292\
        );

    \I__1421\ : InMux
    port map (
            O => \N__6339\,
            I => \N__6292\
        );

    \I__1420\ : InMux
    port map (
            O => \N__6338\,
            I => \N__6292\
        );

    \I__1419\ : InMux
    port map (
            O => \N__6337\,
            I => \N__6286\
        );

    \I__1418\ : InMux
    port map (
            O => \N__6336\,
            I => \N__6286\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__6333\,
            I => \N__6277\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__6324\,
            I => \N__6277\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__6319\,
            I => \N__6277\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__6314\,
            I => \N__6277\
        );

    \I__1413\ : InMux
    port map (
            O => \N__6313\,
            I => \N__6266\
        );

    \I__1412\ : InMux
    port map (
            O => \N__6312\,
            I => \N__6266\
        );

    \I__1411\ : InMux
    port map (
            O => \N__6311\,
            I => \N__6266\
        );

    \I__1410\ : InMux
    port map (
            O => \N__6310\,
            I => \N__6266\
        );

    \I__1409\ : InMux
    port map (
            O => \N__6309\,
            I => \N__6266\
        );

    \I__1408\ : InMux
    port map (
            O => \N__6308\,
            I => \N__6259\
        );

    \I__1407\ : InMux
    port map (
            O => \N__6307\,
            I => \N__6259\
        );

    \I__1406\ : InMux
    port map (
            O => \N__6306\,
            I => \N__6259\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__6301\,
            I => \N__6256\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__6292\,
            I => \N__6253\
        );

    \I__1403\ : InMux
    port map (
            O => \N__6291\,
            I => \N__6250\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__6286\,
            I => \N__6239\
        );

    \I__1401\ : Span4Mux_s3_v
    port map (
            O => \N__6277\,
            I => \N__6239\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__6266\,
            I => \N__6239\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__6259\,
            I => \N__6236\
        );

    \I__1398\ : Span4Mux_s1_v
    port map (
            O => \N__6256\,
            I => \N__6229\
        );

    \I__1397\ : Span4Mux_h
    port map (
            O => \N__6253\,
            I => \N__6229\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__6250\,
            I => \N__6229\
        );

    \I__1395\ : InMux
    port map (
            O => \N__6249\,
            I => \N__6226\
        );

    \I__1394\ : InMux
    port map (
            O => \N__6248\,
            I => \N__6223\
        );

    \I__1393\ : InMux
    port map (
            O => \N__6247\,
            I => \N__6218\
        );

    \I__1392\ : InMux
    port map (
            O => \N__6246\,
            I => \N__6218\
        );

    \I__1391\ : Span4Mux_h
    port map (
            O => \N__6239\,
            I => \N__6215\
        );

    \I__1390\ : Odrv12
    port map (
            O => \N__6236\,
            I => \Gl_rst\
        );

    \I__1389\ : Odrv4
    port map (
            O => \N__6229\,
            I => \Gl_rst\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__6226\,
            I => \Gl_rst\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__6223\,
            I => \Gl_rst\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__6218\,
            I => \Gl_rst\
        );

    \I__1385\ : Odrv4
    port map (
            O => \N__6215\,
            I => \Gl_rst\
        );

    \I__1384\ : InMux
    port map (
            O => \N__6202\,
            I => \N__6199\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__6199\,
            I => \N__6196\
        );

    \I__1382\ : Odrv4
    port map (
            O => \N__6196\,
            I => \L2_adder_rdy\
        );

    \I__1381\ : ClkMux
    port map (
            O => \N__6193\,
            I => \N__6097\
        );

    \I__1380\ : ClkMux
    port map (
            O => \N__6192\,
            I => \N__6097\
        );

    \I__1379\ : ClkMux
    port map (
            O => \N__6191\,
            I => \N__6097\
        );

    \I__1378\ : ClkMux
    port map (
            O => \N__6190\,
            I => \N__6097\
        );

    \I__1377\ : ClkMux
    port map (
            O => \N__6189\,
            I => \N__6097\
        );

    \I__1376\ : ClkMux
    port map (
            O => \N__6188\,
            I => \N__6097\
        );

    \I__1375\ : ClkMux
    port map (
            O => \N__6187\,
            I => \N__6097\
        );

    \I__1374\ : ClkMux
    port map (
            O => \N__6186\,
            I => \N__6097\
        );

    \I__1373\ : ClkMux
    port map (
            O => \N__6185\,
            I => \N__6097\
        );

    \I__1372\ : ClkMux
    port map (
            O => \N__6184\,
            I => \N__6097\
        );

    \I__1371\ : ClkMux
    port map (
            O => \N__6183\,
            I => \N__6097\
        );

    \I__1370\ : ClkMux
    port map (
            O => \N__6182\,
            I => \N__6097\
        );

    \I__1369\ : ClkMux
    port map (
            O => \N__6181\,
            I => \N__6097\
        );

    \I__1368\ : ClkMux
    port map (
            O => \N__6180\,
            I => \N__6097\
        );

    \I__1367\ : ClkMux
    port map (
            O => \N__6179\,
            I => \N__6097\
        );

    \I__1366\ : ClkMux
    port map (
            O => \N__6178\,
            I => \N__6097\
        );

    \I__1365\ : ClkMux
    port map (
            O => \N__6177\,
            I => \N__6097\
        );

    \I__1364\ : ClkMux
    port map (
            O => \N__6176\,
            I => \N__6097\
        );

    \I__1363\ : ClkMux
    port map (
            O => \N__6175\,
            I => \N__6097\
        );

    \I__1362\ : ClkMux
    port map (
            O => \N__6174\,
            I => \N__6097\
        );

    \I__1361\ : ClkMux
    port map (
            O => \N__6173\,
            I => \N__6097\
        );

    \I__1360\ : ClkMux
    port map (
            O => \N__6172\,
            I => \N__6097\
        );

    \I__1359\ : ClkMux
    port map (
            O => \N__6171\,
            I => \N__6097\
        );

    \I__1358\ : ClkMux
    port map (
            O => \N__6170\,
            I => \N__6097\
        );

    \I__1357\ : ClkMux
    port map (
            O => \N__6169\,
            I => \N__6097\
        );

    \I__1356\ : ClkMux
    port map (
            O => \N__6168\,
            I => \N__6097\
        );

    \I__1355\ : ClkMux
    port map (
            O => \N__6167\,
            I => \N__6097\
        );

    \I__1354\ : ClkMux
    port map (
            O => \N__6166\,
            I => \N__6097\
        );

    \I__1353\ : ClkMux
    port map (
            O => \N__6165\,
            I => \N__6097\
        );

    \I__1352\ : ClkMux
    port map (
            O => \N__6164\,
            I => \N__6097\
        );

    \I__1351\ : ClkMux
    port map (
            O => \N__6163\,
            I => \N__6097\
        );

    \I__1350\ : ClkMux
    port map (
            O => \N__6162\,
            I => \N__6097\
        );

    \I__1349\ : GlobalMux
    port map (
            O => \N__6097\,
            I => \N__6094\
        );

    \I__1348\ : gio2CtrlBuf
    port map (
            O => \N__6094\,
            I => clk_g
        );

    \I__1347\ : InMux
    port map (
            O => \N__6091\,
            I => \N__6087\
        );

    \I__1346\ : InMux
    port map (
            O => \N__6090\,
            I => \N__6084\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__6087\,
            I => \N__6081\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__6084\,
            I => \N__6076\
        );

    \I__1343\ : Span4Mux_v
    port map (
            O => \N__6081\,
            I => \N__6076\
        );

    \I__1342\ : Odrv4
    port map (
            O => \N__6076\,
            I => \buart__rx_shifter_fast_4\
        );

    \I__1341\ : CEMux
    port map (
            O => \N__6073\,
            I => \N__6068\
        );

    \I__1340\ : CEMux
    port map (
            O => \N__6072\,
            I => \N__6065\
        );

    \I__1339\ : CEMux
    port map (
            O => \N__6071\,
            I => \N__6062\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__6068\,
            I => \N__6059\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__6065\,
            I => \N__6055\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__6062\,
            I => \N__6052\
        );

    \I__1335\ : Span4Mux_v
    port map (
            O => \N__6059\,
            I => \N__6049\
        );

    \I__1334\ : CEMux
    port map (
            O => \N__6058\,
            I => \N__6046\
        );

    \I__1333\ : Span4Mux_v
    port map (
            O => \N__6055\,
            I => \N__6041\
        );

    \I__1332\ : Span4Mux_s1_h
    port map (
            O => \N__6052\,
            I => \N__6041\
        );

    \I__1331\ : Span4Mux_s2_v
    port map (
            O => \N__6049\,
            I => \N__6036\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__6046\,
            I => \N__6036\
        );

    \I__1329\ : Odrv4
    port map (
            O => \N__6041\,
            I => \buart.Z_rx.sample\
        );

    \I__1328\ : Odrv4
    port map (
            O => \N__6036\,
            I => \buart.Z_rx.sample\
        );

    \I__1327\ : InMux
    port map (
            O => \N__6031\,
            I => \N__6026\
        );

    \I__1326\ : InMux
    port map (
            O => \N__6030\,
            I => \N__6020\
        );

    \I__1325\ : InMux
    port map (
            O => \N__6029\,
            I => \N__6020\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__6026\,
            I => \N__6017\
        );

    \I__1323\ : InMux
    port map (
            O => \N__6025\,
            I => \N__6014\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__6020\,
            I => \Glue_Lab2_Gl_Op_0\
        );

    \I__1321\ : Odrv12
    port map (
            O => \N__6017\,
            I => \Glue_Lab2_Gl_Op_0\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__6014\,
            I => \Glue_Lab2_Gl_Op_0\
        );

    \I__1319\ : InMux
    port map (
            O => \N__6007\,
            I => \N__6002\
        );

    \I__1318\ : InMux
    port map (
            O => \N__6006\,
            I => \N__5996\
        );

    \I__1317\ : InMux
    port map (
            O => \N__6005\,
            I => \N__5996\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__6002\,
            I => \N__5993\
        );

    \I__1315\ : InMux
    port map (
            O => \N__6001\,
            I => \N__5990\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__5996\,
            I => \Glue_Lab2_Gl_Op_3\
        );

    \I__1313\ : Odrv4
    port map (
            O => \N__5993\,
            I => \Glue_Lab2_Gl_Op_3\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__5990\,
            I => \Glue_Lab2_Gl_Op_3\
        );

    \I__1311\ : InMux
    port map (
            O => \N__5983\,
            I => \N__5978\
        );

    \I__1310\ : CascadeMux
    port map (
            O => \N__5982\,
            I => \N__5974\
        );

    \I__1309\ : InMux
    port map (
            O => \N__5981\,
            I => \N__5971\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__5978\,
            I => \N__5968\
        );

    \I__1307\ : InMux
    port map (
            O => \N__5977\,
            I => \N__5963\
        );

    \I__1306\ : InMux
    port map (
            O => \N__5974\,
            I => \N__5963\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__5971\,
            I => \N__5960\
        );

    \I__1304\ : Odrv4
    port map (
            O => \N__5968\,
            I => \Glue_Lab2_Gl_Op_1\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__5963\,
            I => \Glue_Lab2_Gl_Op_1\
        );

    \I__1302\ : Odrv4
    port map (
            O => \N__5960\,
            I => \Glue_Lab2_Gl_Op_1\
        );

    \I__1301\ : InMux
    port map (
            O => \N__5953\,
            I => \N__5947\
        );

    \I__1300\ : InMux
    port map (
            O => \N__5952\,
            I => \N__5944\
        );

    \I__1299\ : InMux
    port map (
            O => \N__5951\,
            I => \N__5941\
        );

    \I__1298\ : InMux
    port map (
            O => \N__5950\,
            I => \N__5938\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__5947\,
            I => \N__5935\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__5944\,
            I => \N__5932\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__5941\,
            I => \Glue_Lab2_Gl_Op_5\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__5938\,
            I => \Glue_Lab2_Gl_Op_5\
        );

    \I__1293\ : Odrv4
    port map (
            O => \N__5935\,
            I => \Glue_Lab2_Gl_Op_5\
        );

    \I__1292\ : Odrv4
    port map (
            O => \N__5932\,
            I => \Glue_Lab2_Gl_Op_5\
        );

    \I__1291\ : CascadeMux
    port map (
            O => \N__5923\,
            I => \Glue_Lab2.g0_0_1_0_cascade_\
        );

    \I__1290\ : InMux
    port map (
            O => \N__5920\,
            I => \N__5917\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__5917\,
            I => \N__5911\
        );

    \I__1288\ : InMux
    port map (
            O => \N__5916\,
            I => \N__5906\
        );

    \I__1287\ : InMux
    port map (
            O => \N__5915\,
            I => \N__5906\
        );

    \I__1286\ : InMux
    port map (
            O => \N__5914\,
            I => \N__5903\
        );

    \I__1285\ : Odrv12
    port map (
            O => \N__5911\,
            I => \Glue_Lab2_Gl_Op_2\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__5906\,
            I => \Glue_Lab2_Gl_Op_2\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__5903\,
            I => \Glue_Lab2_Gl_Op_2\
        );

    \I__1282\ : InMux
    port map (
            O => \N__5896\,
            I => \N__5893\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__5893\,
            I => \N__5890\
        );

    \I__1280\ : Span4Mux_h
    port map (
            O => \N__5890\,
            I => \N__5887\
        );

    \I__1279\ : Odrv4
    port map (
            O => \N__5887\,
            I => \Glue_Lab2.Gl_subtract_0\
        );

    \I__1278\ : InMux
    port map (
            O => \N__5884\,
            I => \N__5877\
        );

    \I__1277\ : InMux
    port map (
            O => \N__5883\,
            I => \N__5877\
        );

    \I__1276\ : InMux
    port map (
            O => \N__5882\,
            I => \N__5874\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__5877\,
            I => \N__5868\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__5874\,
            I => \N__5865\
        );

    \I__1273\ : InMux
    port map (
            O => \N__5873\,
            I => \N__5857\
        );

    \I__1272\ : InMux
    port map (
            O => \N__5872\,
            I => \N__5854\
        );

    \I__1271\ : InMux
    port map (
            O => \N__5871\,
            I => \N__5851\
        );

    \I__1270\ : Span4Mux_h
    port map (
            O => \N__5868\,
            I => \N__5846\
        );

    \I__1269\ : Span4Mux_h
    port map (
            O => \N__5865\,
            I => \N__5846\
        );

    \I__1268\ : InMux
    port map (
            O => \N__5864\,
            I => \N__5841\
        );

    \I__1267\ : InMux
    port map (
            O => \N__5863\,
            I => \N__5841\
        );

    \I__1266\ : InMux
    port map (
            O => \N__5862\,
            I => \N__5836\
        );

    \I__1265\ : InMux
    port map (
            O => \N__5861\,
            I => \N__5836\
        );

    \I__1264\ : InMux
    port map (
            O => \N__5860\,
            I => \N__5833\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__5857\,
            I => \N__5830\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__5854\,
            I => \Gl_r1_2\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__5851\,
            I => \Gl_r1_2\
        );

    \I__1260\ : Odrv4
    port map (
            O => \N__5846\,
            I => \Gl_r1_2\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__5841\,
            I => \Gl_r1_2\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__5836\,
            I => \Gl_r1_2\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__5833\,
            I => \Gl_r1_2\
        );

    \I__1256\ : Odrv4
    port map (
            O => \N__5830\,
            I => \Gl_r1_2\
        );

    \I__1255\ : InMux
    port map (
            O => \N__5815\,
            I => \N__5806\
        );

    \I__1254\ : InMux
    port map (
            O => \N__5814\,
            I => \N__5806\
        );

    \I__1253\ : InMux
    port map (
            O => \N__5813\,
            I => \N__5802\
        );

    \I__1252\ : CascadeMux
    port map (
            O => \N__5812\,
            I => \N__5797\
        );

    \I__1251\ : CascadeMux
    port map (
            O => \N__5811\,
            I => \N__5794\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__5806\,
            I => \N__5791\
        );

    \I__1249\ : InMux
    port map (
            O => \N__5805\,
            I => \N__5788\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__5802\,
            I => \N__5785\
        );

    \I__1247\ : CascadeMux
    port map (
            O => \N__5801\,
            I => \N__5781\
        );

    \I__1246\ : InMux
    port map (
            O => \N__5800\,
            I => \N__5776\
        );

    \I__1245\ : InMux
    port map (
            O => \N__5797\,
            I => \N__5773\
        );

    \I__1244\ : InMux
    port map (
            O => \N__5794\,
            I => \N__5770\
        );

    \I__1243\ : Span4Mux_h
    port map (
            O => \N__5791\,
            I => \N__5763\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__5788\,
            I => \N__5763\
        );

    \I__1241\ : Span4Mux_h
    port map (
            O => \N__5785\,
            I => \N__5763\
        );

    \I__1240\ : InMux
    port map (
            O => \N__5784\,
            I => \N__5760\
        );

    \I__1239\ : InMux
    port map (
            O => \N__5781\,
            I => \N__5757\
        );

    \I__1238\ : InMux
    port map (
            O => \N__5780\,
            I => \N__5752\
        );

    \I__1237\ : InMux
    port map (
            O => \N__5779\,
            I => \N__5752\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__5776\,
            I => \N__5749\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__5773\,
            I => \Gl_r2_2\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__5770\,
            I => \Gl_r2_2\
        );

    \I__1233\ : Odrv4
    port map (
            O => \N__5763\,
            I => \Gl_r2_2\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__5760\,
            I => \Gl_r2_2\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__5757\,
            I => \Gl_r2_2\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__5752\,
            I => \Gl_r2_2\
        );

    \I__1229\ : Odrv4
    port map (
            O => \N__5749\,
            I => \Gl_r2_2\
        );

    \I__1228\ : InMux
    port map (
            O => \N__5734\,
            I => \N__5728\
        );

    \I__1227\ : InMux
    port map (
            O => \N__5733\,
            I => \N__5728\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__5728\,
            I => \N__5725\
        );

    \I__1225\ : Span4Mux_h
    port map (
            O => \N__5725\,
            I => \N__5712\
        );

    \I__1224\ : InMux
    port map (
            O => \N__5724\,
            I => \N__5707\
        );

    \I__1223\ : InMux
    port map (
            O => \N__5723\,
            I => \N__5707\
        );

    \I__1222\ : InMux
    port map (
            O => \N__5722\,
            I => \N__5702\
        );

    \I__1221\ : InMux
    port map (
            O => \N__5721\,
            I => \N__5702\
        );

    \I__1220\ : InMux
    port map (
            O => \N__5720\,
            I => \N__5695\
        );

    \I__1219\ : InMux
    port map (
            O => \N__5719\,
            I => \N__5695\
        );

    \I__1218\ : InMux
    port map (
            O => \N__5718\,
            I => \N__5695\
        );

    \I__1217\ : InMux
    port map (
            O => \N__5717\,
            I => \N__5688\
        );

    \I__1216\ : InMux
    port map (
            O => \N__5716\,
            I => \N__5688\
        );

    \I__1215\ : InMux
    port map (
            O => \N__5715\,
            I => \N__5688\
        );

    \I__1214\ : Odrv4
    port map (
            O => \N__5712\,
            I => \Gl_r1_3\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__5707\,
            I => \Gl_r1_3\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__5702\,
            I => \Gl_r1_3\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__5695\,
            I => \Gl_r1_3\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__5688\,
            I => \Gl_r1_3\
        );

    \I__1209\ : InMux
    port map (
            O => \N__5677\,
            I => \N__5674\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__5674\,
            I => \N__5671\
        );

    \I__1207\ : Span4Mux_v
    port map (
            O => \N__5671\,
            I => \N__5668\
        );

    \I__1206\ : Odrv4
    port map (
            O => \N__5668\,
            I => \Lab_UT.S_1_c3_d\
        );

    \I__1205\ : CascadeMux
    port map (
            O => \N__5665\,
            I => \Lab_UT.S_1_c3_cZ0_cascade_\
        );

    \I__1204\ : CascadeMux
    port map (
            O => \N__5662\,
            I => \N__5657\
        );

    \I__1203\ : CascadeMux
    port map (
            O => \N__5661\,
            I => \N__5653\
        );

    \I__1202\ : InMux
    port map (
            O => \N__5660\,
            I => \N__5646\
        );

    \I__1201\ : InMux
    port map (
            O => \N__5657\,
            I => \N__5646\
        );

    \I__1200\ : CascadeMux
    port map (
            O => \N__5656\,
            I => \N__5643\
        );

    \I__1199\ : InMux
    port map (
            O => \N__5653\,
            I => \N__5634\
        );

    \I__1198\ : InMux
    port map (
            O => \N__5652\,
            I => \N__5634\
        );

    \I__1197\ : InMux
    port map (
            O => \N__5651\,
            I => \N__5634\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__5646\,
            I => \N__5627\
        );

    \I__1195\ : InMux
    port map (
            O => \N__5643\,
            I => \N__5620\
        );

    \I__1194\ : InMux
    port map (
            O => \N__5642\,
            I => \N__5620\
        );

    \I__1193\ : InMux
    port map (
            O => \N__5641\,
            I => \N__5620\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__5634\,
            I => \N__5617\
        );

    \I__1191\ : InMux
    port map (
            O => \N__5633\,
            I => \N__5612\
        );

    \I__1190\ : InMux
    port map (
            O => \N__5632\,
            I => \N__5612\
        );

    \I__1189\ : InMux
    port map (
            O => \N__5631\,
            I => \N__5607\
        );

    \I__1188\ : InMux
    port map (
            O => \N__5630\,
            I => \N__5607\
        );

    \I__1187\ : Span4Mux_h
    port map (
            O => \N__5627\,
            I => \N__5602\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__5620\,
            I => \N__5602\
        );

    \I__1185\ : Odrv4
    port map (
            O => \N__5617\,
            I => \Gl_r2_3\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__5612\,
            I => \Gl_r2_3\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__5607\,
            I => \Gl_r2_3\
        );

    \I__1182\ : Odrv4
    port map (
            O => \N__5602\,
            I => \Gl_r2_3\
        );

    \I__1181\ : InMux
    port map (
            O => \N__5593\,
            I => \N__5590\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__5590\,
            I => \Lab_UT.S_0_s_ac0_5_0Z0Z_0\
        );

    \I__1179\ : InMux
    port map (
            O => \N__5587\,
            I => \N__5584\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__5584\,
            I => \N__5581\
        );

    \I__1177\ : Span4Mux_v
    port map (
            O => \N__5581\,
            I => \N__5578\
        );

    \I__1176\ : Odrv4
    port map (
            O => \N__5578\,
            I => \Lab_UT.S_0_s_ac0_5_dZ0\
        );

    \I__1175\ : CascadeMux
    port map (
            O => \N__5575\,
            I => \Lab_UT.C_out41_cascade_\
        );

    \I__1174\ : InMux
    port map (
            O => \N__5572\,
            I => \N__5568\
        );

    \I__1173\ : InMux
    port map (
            O => \N__5571\,
            I => \N__5565\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__5568\,
            I => \N__5562\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__5565\,
            I => \N__5559\
        );

    \I__1170\ : Span4Mux_s3_h
    port map (
            O => \N__5562\,
            I => \N__5552\
        );

    \I__1169\ : Span4Mux_h
    port map (
            O => \N__5559\,
            I => \N__5552\
        );

    \I__1168\ : InMux
    port map (
            O => \N__5558\,
            I => \N__5547\
        );

    \I__1167\ : InMux
    port map (
            O => \N__5557\,
            I => \N__5547\
        );

    \I__1166\ : Odrv4
    port map (
            O => \N__5552\,
            I => \Gl_subtract\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__5547\,
            I => \Gl_subtract\
        );

    \I__1164\ : IoInMux
    port map (
            O => \N__5542\,
            I => \N__5539\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__5539\,
            I => \N__5536\
        );

    \I__1162\ : Span4Mux_s2_h
    port map (
            O => \N__5536\,
            I => \N__5533\
        );

    \I__1161\ : Span4Mux_v
    port map (
            O => \N__5533\,
            I => \N__5530\
        );

    \I__1160\ : Odrv4
    port map (
            O => \N__5530\,
            I => led_c_4
        );

    \I__1159\ : CascadeMux
    port map (
            O => \N__5527\,
            I => \Glue_Lab2.de0.g0_5_1_cascade_\
        );

    \I__1158\ : CascadeMux
    port map (
            O => \N__5524\,
            I => \Glue_Lab2.g0_9_1_cascade_\
        );

    \I__1157\ : InMux
    port map (
            O => \N__5521\,
            I => \N__5518\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__5518\,
            I => \N__5515\
        );

    \I__1155\ : Span4Mux_v
    port map (
            O => \N__5515\,
            I => \N__5512\
        );

    \I__1154\ : Odrv4
    port map (
            O => \N__5512\,
            I => \Glue_Lab2.g0_7_1\
        );

    \I__1153\ : InMux
    port map (
            O => \N__5509\,
            I => \N__5506\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__5506\,
            I => \N__5503\
        );

    \I__1151\ : Odrv12
    port map (
            O => \N__5503\,
            I => \Glue_Lab2.reset_counte_0_2\
        );

    \I__1150\ : InMux
    port map (
            O => \N__5500\,
            I => \N__5496\
        );

    \I__1149\ : InMux
    port map (
            O => \N__5499\,
            I => \N__5490\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__5496\,
            I => \N__5484\
        );

    \I__1147\ : InMux
    port map (
            O => \N__5495\,
            I => \N__5477\
        );

    \I__1146\ : InMux
    port map (
            O => \N__5494\,
            I => \N__5477\
        );

    \I__1145\ : InMux
    port map (
            O => \N__5493\,
            I => \N__5477\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__5490\,
            I => \N__5474\
        );

    \I__1143\ : InMux
    port map (
            O => \N__5489\,
            I => \N__5467\
        );

    \I__1142\ : InMux
    port map (
            O => \N__5488\,
            I => \N__5467\
        );

    \I__1141\ : InMux
    port map (
            O => \N__5487\,
            I => \N__5467\
        );

    \I__1140\ : Span4Mux_v
    port map (
            O => \N__5484\,
            I => \N__5462\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__5477\,
            I => \N__5462\
        );

    \I__1138\ : Odrv4
    port map (
            O => \N__5474\,
            I => bu_rx_data_4
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__5467\,
            I => bu_rx_data_4
        );

    \I__1136\ : Odrv4
    port map (
            O => \N__5462\,
            I => bu_rx_data_4
        );

    \I__1135\ : InMux
    port map (
            O => \N__5455\,
            I => \N__5448\
        );

    \I__1134\ : InMux
    port map (
            O => \N__5454\,
            I => \N__5448\
        );

    \I__1133\ : InMux
    port map (
            O => \N__5453\,
            I => \N__5444\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__5448\,
            I => \N__5440\
        );

    \I__1131\ : InMux
    port map (
            O => \N__5447\,
            I => \N__5432\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__5444\,
            I => \N__5429\
        );

    \I__1129\ : InMux
    port map (
            O => \N__5443\,
            I => \N__5426\
        );

    \I__1128\ : Span4Mux_s3_h
    port map (
            O => \N__5440\,
            I => \N__5423\
        );

    \I__1127\ : InMux
    port map (
            O => \N__5439\,
            I => \N__5420\
        );

    \I__1126\ : InMux
    port map (
            O => \N__5438\,
            I => \N__5417\
        );

    \I__1125\ : InMux
    port map (
            O => \N__5437\,
            I => \N__5414\
        );

    \I__1124\ : InMux
    port map (
            O => \N__5436\,
            I => \N__5409\
        );

    \I__1123\ : InMux
    port map (
            O => \N__5435\,
            I => \N__5409\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__5432\,
            I => \buart__rx_bitcount_0\
        );

    \I__1121\ : Odrv4
    port map (
            O => \N__5429\,
            I => \buart__rx_bitcount_0\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__5426\,
            I => \buart__rx_bitcount_0\
        );

    \I__1119\ : Odrv4
    port map (
            O => \N__5423\,
            I => \buart__rx_bitcount_0\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__5420\,
            I => \buart__rx_bitcount_0\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__5417\,
            I => \buart__rx_bitcount_0\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__5414\,
            I => \buart__rx_bitcount_0\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__5409\,
            I => \buart__rx_bitcount_0\
        );

    \I__1114\ : CascadeMux
    port map (
            O => \N__5392\,
            I => \Glue_Lab2.de0.g0Z0Z_5_cascade_\
        );

    \I__1113\ : InMux
    port map (
            O => \N__5389\,
            I => \N__5377\
        );

    \I__1112\ : InMux
    port map (
            O => \N__5388\,
            I => \N__5377\
        );

    \I__1111\ : InMux
    port map (
            O => \N__5387\,
            I => \N__5374\
        );

    \I__1110\ : InMux
    port map (
            O => \N__5386\,
            I => \N__5371\
        );

    \I__1109\ : InMux
    port map (
            O => \N__5385\,
            I => \N__5366\
        );

    \I__1108\ : InMux
    port map (
            O => \N__5384\,
            I => \N__5366\
        );

    \I__1107\ : InMux
    port map (
            O => \N__5383\,
            I => \N__5363\
        );

    \I__1106\ : InMux
    port map (
            O => \N__5382\,
            I => \N__5360\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__5377\,
            I => \N__5357\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__5374\,
            I => \N__5352\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__5371\,
            I => \N__5349\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__5366\,
            I => \N__5346\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__5363\,
            I => \N__5341\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__5360\,
            I => \N__5336\
        );

    \I__1099\ : Span4Mux_v
    port map (
            O => \N__5357\,
            I => \N__5336\
        );

    \I__1098\ : InMux
    port map (
            O => \N__5356\,
            I => \N__5331\
        );

    \I__1097\ : InMux
    port map (
            O => \N__5355\,
            I => \N__5331\
        );

    \I__1096\ : Span4Mux_h
    port map (
            O => \N__5352\,
            I => \N__5328\
        );

    \I__1095\ : Span4Mux_h
    port map (
            O => \N__5349\,
            I => \N__5323\
        );

    \I__1094\ : Span4Mux_s2_h
    port map (
            O => \N__5346\,
            I => \N__5323\
        );

    \I__1093\ : InMux
    port map (
            O => \N__5345\,
            I => \N__5318\
        );

    \I__1092\ : InMux
    port map (
            O => \N__5344\,
            I => \N__5318\
        );

    \I__1091\ : Odrv4
    port map (
            O => \N__5341\,
            I => bu_rx_data_0
        );

    \I__1090\ : Odrv4
    port map (
            O => \N__5336\,
            I => bu_rx_data_0
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__5331\,
            I => bu_rx_data_0
        );

    \I__1088\ : Odrv4
    port map (
            O => \N__5328\,
            I => bu_rx_data_0
        );

    \I__1087\ : Odrv4
    port map (
            O => \N__5323\,
            I => bu_rx_data_0
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__5318\,
            I => bu_rx_data_0
        );

    \I__1085\ : InMux
    port map (
            O => \N__5305\,
            I => \N__5300\
        );

    \I__1084\ : InMux
    port map (
            O => \N__5304\,
            I => \N__5295\
        );

    \I__1083\ : InMux
    port map (
            O => \N__5303\,
            I => \N__5295\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__5300\,
            I => \N__5289\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__5295\,
            I => \N__5286\
        );

    \I__1080\ : InMux
    port map (
            O => \N__5294\,
            I => \N__5283\
        );

    \I__1079\ : InMux
    port map (
            O => \N__5293\,
            I => \N__5280\
        );

    \I__1078\ : InMux
    port map (
            O => \N__5292\,
            I => \N__5277\
        );

    \I__1077\ : Span4Mux_h
    port map (
            O => \N__5289\,
            I => \N__5274\
        );

    \I__1076\ : Span4Mux_s2_h
    port map (
            O => \N__5286\,
            I => \N__5269\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__5283\,
            I => \N__5269\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__5280\,
            I => \Glue_Lab2.reset_countZ0Z_4\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__5277\,
            I => \Glue_Lab2.reset_countZ0Z_4\
        );

    \I__1072\ : Odrv4
    port map (
            O => \N__5274\,
            I => \Glue_Lab2.reset_countZ0Z_4\
        );

    \I__1071\ : Odrv4
    port map (
            O => \N__5269\,
            I => \Glue_Lab2.reset_countZ0Z_4\
        );

    \I__1070\ : CascadeMux
    port map (
            O => \N__5260\,
            I => \Glue_Lab2.g0_9_cascade_\
        );

    \I__1069\ : InMux
    port map (
            O => \N__5257\,
            I => \N__5254\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__5254\,
            I => \N__5251\
        );

    \I__1067\ : Odrv4
    port map (
            O => \N__5251\,
            I => \Glue_Lab2.g0_7\
        );

    \I__1066\ : InMux
    port map (
            O => \N__5248\,
            I => \N__5245\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__5245\,
            I => \N__5242\
        );

    \I__1064\ : Span4Mux_h
    port map (
            O => \N__5242\,
            I => \N__5239\
        );

    \I__1063\ : Odrv4
    port map (
            O => \N__5239\,
            I => \Glue_Lab2.reset_counte_0_0\
        );

    \I__1062\ : InMux
    port map (
            O => \N__5236\,
            I => \N__5223\
        );

    \I__1061\ : InMux
    port map (
            O => \N__5235\,
            I => \N__5220\
        );

    \I__1060\ : InMux
    port map (
            O => \N__5234\,
            I => \N__5213\
        );

    \I__1059\ : InMux
    port map (
            O => \N__5233\,
            I => \N__5213\
        );

    \I__1058\ : InMux
    port map (
            O => \N__5232\,
            I => \N__5213\
        );

    \I__1057\ : InMux
    port map (
            O => \N__5231\,
            I => \N__5210\
        );

    \I__1056\ : InMux
    port map (
            O => \N__5230\,
            I => \N__5207\
        );

    \I__1055\ : InMux
    port map (
            O => \N__5229\,
            I => \N__5204\
        );

    \I__1054\ : InMux
    port map (
            O => \N__5228\,
            I => \N__5201\
        );

    \I__1053\ : InMux
    port map (
            O => \N__5227\,
            I => \N__5198\
        );

    \I__1052\ : InMux
    port map (
            O => \N__5226\,
            I => \N__5193\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__5223\,
            I => \N__5184\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__5220\,
            I => \N__5184\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__5213\,
            I => \N__5184\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__5210\,
            I => \N__5184\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__5207\,
            I => \N__5181\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__5204\,
            I => \N__5178\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__5201\,
            I => \N__5170\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__5198\,
            I => \N__5170\
        );

    \I__1043\ : InMux
    port map (
            O => \N__5197\,
            I => \N__5167\
        );

    \I__1042\ : InMux
    port map (
            O => \N__5196\,
            I => \N__5164\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__5193\,
            I => \N__5157\
        );

    \I__1040\ : Span4Mux_v
    port map (
            O => \N__5184\,
            I => \N__5157\
        );

    \I__1039\ : Span4Mux_v
    port map (
            O => \N__5181\,
            I => \N__5157\
        );

    \I__1038\ : Span4Mux_h
    port map (
            O => \N__5178\,
            I => \N__5154\
        );

    \I__1037\ : InMux
    port map (
            O => \N__5177\,
            I => \N__5147\
        );

    \I__1036\ : InMux
    port map (
            O => \N__5176\,
            I => \N__5147\
        );

    \I__1035\ : InMux
    port map (
            O => \N__5175\,
            I => \N__5147\
        );

    \I__1034\ : Span12Mux_s4_v
    port map (
            O => \N__5170\,
            I => \N__5140\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__5167\,
            I => \N__5140\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__5164\,
            I => \N__5140\
        );

    \I__1031\ : Odrv4
    port map (
            O => \N__5157\,
            I => bu_rx_data_2
        );

    \I__1030\ : Odrv4
    port map (
            O => \N__5154\,
            I => bu_rx_data_2
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__5147\,
            I => bu_rx_data_2
        );

    \I__1028\ : Odrv12
    port map (
            O => \N__5140\,
            I => bu_rx_data_2
        );

    \I__1027\ : InMux
    port map (
            O => \N__5131\,
            I => \N__5126\
        );

    \I__1026\ : InMux
    port map (
            O => \N__5130\,
            I => \N__5123\
        );

    \I__1025\ : CascadeMux
    port map (
            O => \N__5129\,
            I => \N__5120\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__5126\,
            I => \N__5115\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__5123\,
            I => \N__5112\
        );

    \I__1022\ : InMux
    port map (
            O => \N__5120\,
            I => \N__5105\
        );

    \I__1021\ : InMux
    port map (
            O => \N__5119\,
            I => \N__5105\
        );

    \I__1020\ : InMux
    port map (
            O => \N__5118\,
            I => \N__5105\
        );

    \I__1019\ : Span4Mux_v
    port map (
            O => \N__5115\,
            I => \N__5092\
        );

    \I__1018\ : Span4Mux_v
    port map (
            O => \N__5112\,
            I => \N__5092\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__5105\,
            I => \N__5092\
        );

    \I__1016\ : InMux
    port map (
            O => \N__5104\,
            I => \N__5089\
        );

    \I__1015\ : InMux
    port map (
            O => \N__5103\,
            I => \N__5080\
        );

    \I__1014\ : InMux
    port map (
            O => \N__5102\,
            I => \N__5080\
        );

    \I__1013\ : InMux
    port map (
            O => \N__5101\,
            I => \N__5080\
        );

    \I__1012\ : InMux
    port map (
            O => \N__5100\,
            I => \N__5080\
        );

    \I__1011\ : InMux
    port map (
            O => \N__5099\,
            I => \N__5077\
        );

    \I__1010\ : Odrv4
    port map (
            O => \N__5092\,
            I => bu_rx_data_6
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__5089\,
            I => bu_rx_data_6
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__5080\,
            I => bu_rx_data_6
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__5077\,
            I => bu_rx_data_6
        );

    \I__1006\ : InMux
    port map (
            O => \N__5068\,
            I => \N__5059\
        );

    \I__1005\ : InMux
    port map (
            O => \N__5067\,
            I => \N__5059\
        );

    \I__1004\ : InMux
    port map (
            O => \N__5066\,
            I => \N__5059\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__5059\,
            I => \buart.Z_tx.bitcountZ0Z_2\
        );

    \I__1002\ : CascadeMux
    port map (
            O => \N__5056\,
            I => \buart.Z_tx.un1_bitcount_c3_cascade_\
        );

    \I__1001\ : InMux
    port map (
            O => \N__5053\,
            I => \N__5047\
        );

    \I__1000\ : InMux
    port map (
            O => \N__5052\,
            I => \N__5047\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__5047\,
            I => \buart.Z_tx.bitcountZ0Z_3\
        );

    \I__998\ : InMux
    port map (
            O => \N__5044\,
            I => \N__5041\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__5041\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i_sx\
        );

    \I__996\ : InMux
    port map (
            O => \N__5038\,
            I => \N__5034\
        );

    \I__995\ : CascadeMux
    port map (
            O => \N__5037\,
            I => \N__5028\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__5034\,
            I => \N__5025\
        );

    \I__993\ : InMux
    port map (
            O => \N__5033\,
            I => \N__5022\
        );

    \I__992\ : InMux
    port map (
            O => \N__5032\,
            I => \N__5019\
        );

    \I__991\ : InMux
    port map (
            O => \N__5031\,
            I => \N__5011\
        );

    \I__990\ : InMux
    port map (
            O => \N__5028\,
            I => \N__5011\
        );

    \I__989\ : Span4Mux_s3_h
    port map (
            O => \N__5025\,
            I => \N__5005\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__5022\,
            I => \N__5000\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__5019\,
            I => \N__5000\
        );

    \I__986\ : InMux
    port map (
            O => \N__5018\,
            I => \N__4995\
        );

    \I__985\ : InMux
    port map (
            O => \N__5017\,
            I => \N__4995\
        );

    \I__984\ : InMux
    port map (
            O => \N__5016\,
            I => \N__4992\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__5011\,
            I => \N__4989\
        );

    \I__982\ : InMux
    port map (
            O => \N__5010\,
            I => \N__4982\
        );

    \I__981\ : InMux
    port map (
            O => \N__5009\,
            I => \N__4982\
        );

    \I__980\ : InMux
    port map (
            O => \N__5008\,
            I => \N__4982\
        );

    \I__979\ : Odrv4
    port map (
            O => \N__5005\,
            I => \Glue_Lab2.is_hexplus\
        );

    \I__978\ : Odrv4
    port map (
            O => \N__5000\,
            I => \Glue_Lab2.is_hexplus\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__4995\,
            I => \Glue_Lab2.is_hexplus\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__4992\,
            I => \Glue_Lab2.is_hexplus\
        );

    \I__975\ : Odrv4
    port map (
            O => \N__4989\,
            I => \Glue_Lab2.is_hexplus\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__4982\,
            I => \Glue_Lab2.is_hexplus\
        );

    \I__973\ : CascadeMux
    port map (
            O => \N__4969\,
            I => \buart.Z_tx.un1_bitcount_c1_cascade_\
        );

    \I__972\ : CascadeMux
    port map (
            O => \N__4966\,
            I => \N__4962\
        );

    \I__971\ : InMux
    port map (
            O => \N__4965\,
            I => \N__4956\
        );

    \I__970\ : InMux
    port map (
            O => \N__4962\,
            I => \N__4949\
        );

    \I__969\ : InMux
    port map (
            O => \N__4961\,
            I => \N__4949\
        );

    \I__968\ : InMux
    port map (
            O => \N__4960\,
            I => \N__4949\
        );

    \I__967\ : InMux
    port map (
            O => \N__4959\,
            I => \N__4946\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__4956\,
            I => \buart.Z_tx.bitcountZ0Z_1\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__4949\,
            I => \buart.Z_tx.bitcountZ0Z_1\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__4946\,
            I => \buart.Z_tx.bitcountZ0Z_1\
        );

    \I__963\ : InMux
    port map (
            O => \N__4939\,
            I => \N__4934\
        );

    \I__962\ : InMux
    port map (
            O => \N__4938\,
            I => \N__4929\
        );

    \I__961\ : InMux
    port map (
            O => \N__4937\,
            I => \N__4929\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__4934\,
            I => \buart.Z_tx.counter_RNIVE1P1_4\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__4929\,
            I => \buart.Z_tx.counter_RNIVE1P1_4\
        );

    \I__958\ : InMux
    port map (
            O => \N__4924\,
            I => \N__4914\
        );

    \I__957\ : InMux
    port map (
            O => \N__4923\,
            I => \N__4914\
        );

    \I__956\ : InMux
    port map (
            O => \N__4922\,
            I => \N__4905\
        );

    \I__955\ : InMux
    port map (
            O => \N__4921\,
            I => \N__4905\
        );

    \I__954\ : InMux
    port map (
            O => \N__4920\,
            I => \N__4905\
        );

    \I__953\ : InMux
    port map (
            O => \N__4919\,
            I => \N__4905\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__4914\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__4905\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__950\ : InMux
    port map (
            O => \N__4900\,
            I => \N__4897\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__4897\,
            I => \N__4894\
        );

    \I__948\ : Span4Mux_h
    port map (
            O => \N__4894\,
            I => \N__4891\
        );

    \I__947\ : Odrv4
    port map (
            O => \N__4891\,
            I => \Glue_Lab2.de0.de_escZ0Z_4\
        );

    \I__946\ : InMux
    port map (
            O => \N__4888\,
            I => \N__4876\
        );

    \I__945\ : InMux
    port map (
            O => \N__4887\,
            I => \N__4876\
        );

    \I__944\ : InMux
    port map (
            O => \N__4886\,
            I => \N__4876\
        );

    \I__943\ : InMux
    port map (
            O => \N__4885\,
            I => \N__4876\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__4876\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_4\
        );

    \I__941\ : CascadeMux
    port map (
            O => \N__4873\,
            I => \N__4867\
        );

    \I__940\ : InMux
    port map (
            O => \N__4872\,
            I => \N__4858\
        );

    \I__939\ : InMux
    port map (
            O => \N__4871\,
            I => \N__4858\
        );

    \I__938\ : InMux
    port map (
            O => \N__4870\,
            I => \N__4858\
        );

    \I__937\ : InMux
    port map (
            O => \N__4867\,
            I => \N__4858\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__4858\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_5\
        );

    \I__935\ : InMux
    port map (
            O => \N__4855\,
            I => \N__4846\
        );

    \I__934\ : InMux
    port map (
            O => \N__4854\,
            I => \N__4846\
        );

    \I__933\ : InMux
    port map (
            O => \N__4853\,
            I => \N__4846\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__4846\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_6\
        );

    \I__931\ : CascadeMux
    port map (
            O => \N__4843\,
            I => \N__4840\
        );

    \I__930\ : InMux
    port map (
            O => \N__4840\,
            I => \N__4832\
        );

    \I__929\ : InMux
    port map (
            O => \N__4839\,
            I => \N__4832\
        );

    \I__928\ : InMux
    port map (
            O => \N__4838\,
            I => \N__4827\
        );

    \I__927\ : InMux
    port map (
            O => \N__4837\,
            I => \N__4827\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__4832\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__4827\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__924\ : CascadeMux
    port map (
            O => \N__4822\,
            I => \buart.Z_tx.Z_baudgen.ser_clk_sx_cascade_\
        );

    \I__923\ : InMux
    port map (
            O => \N__4819\,
            I => \N__4808\
        );

    \I__922\ : InMux
    port map (
            O => \N__4818\,
            I => \N__4808\
        );

    \I__921\ : InMux
    port map (
            O => \N__4817\,
            I => \N__4808\
        );

    \I__920\ : InMux
    port map (
            O => \N__4816\,
            I => \N__4803\
        );

    \I__919\ : InMux
    port map (
            O => \N__4815\,
            I => \N__4803\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__4808\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__4803\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__916\ : InMux
    port map (
            O => \N__4798\,
            I => \N__4795\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__4795\,
            I => \buart.Z_tx.Z_baudgen.counter_RNIES38_0Z0Z_4\
        );

    \I__914\ : InMux
    port map (
            O => \N__4792\,
            I => \N__4789\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__4789\,
            I => \buart.Z_tx.Z_baudgen.un1_bitcount_c2_1\
        );

    \I__912\ : CascadeMux
    port map (
            O => \N__4786\,
            I => \buart.Z_tx.bitcount_RNIBADLZ0Z_1_cascade_\
        );

    \I__911\ : CascadeMux
    port map (
            O => \N__4783\,
            I => \buart.Z_tx.counter_RNIVE1P1_4_cascade_\
        );

    \I__910\ : InMux
    port map (
            O => \N__4780\,
            I => \N__4777\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__4777\,
            I => \buart.Z_tx.un1_bitcount_c2\
        );

    \I__908\ : InMux
    port map (
            O => \N__4774\,
            I => \N__4771\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__4771\,
            I => \buart.Z_tx.uart_busy_0_0\
        );

    \I__906\ : CascadeMux
    port map (
            O => \N__4768\,
            I => \buart.Z_tx.uart_busy_0_0_cascade_\
        );

    \I__905\ : CascadeMux
    port map (
            O => \N__4765\,
            I => \led_c_1_cascade_\
        );

    \I__904\ : InMux
    port map (
            O => \N__4762\,
            I => \N__4759\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__4759\,
            I => \N__4756\
        );

    \I__902\ : Span12Mux_s8_h
    port map (
            O => \N__4756\,
            I => \N__4753\
        );

    \I__901\ : Odrv12
    port map (
            O => \N__4753\,
            I => \Gl_tx_data_1\
        );

    \I__900\ : InMux
    port map (
            O => \N__4750\,
            I => \N__4747\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__4747\,
            I => \N__4743\
        );

    \I__898\ : InMux
    port map (
            O => \N__4746\,
            I => \N__4740\
        );

    \I__897\ : Odrv4
    port map (
            O => \N__4743\,
            I => \Gl_r2_fast_2\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__4740\,
            I => \Gl_r2_fast_2\
        );

    \I__895\ : InMux
    port map (
            O => \N__4735\,
            I => \N__4731\
        );

    \I__894\ : InMux
    port map (
            O => \N__4734\,
            I => \N__4728\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__4731\,
            I => \Gl_r1_fast_2\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__4728\,
            I => \Gl_r1_fast_2\
        );

    \I__891\ : InMux
    port map (
            O => \N__4723\,
            I => \N__4720\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__4720\,
            I => \Lab_UT.S_m_bm_1Z0Z_2\
        );

    \I__889\ : InMux
    port map (
            O => \N__4717\,
            I => \N__4714\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__4714\,
            I => \Lab_UT.S_m_bmZ0Z_2\
        );

    \I__887\ : CascadeMux
    port map (
            O => \N__4711\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_c5_cascade_\
        );

    \I__886\ : CascadeMux
    port map (
            O => \N__4708\,
            I => \N__4705\
        );

    \I__885\ : InMux
    port map (
            O => \N__4705\,
            I => \N__4702\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__4702\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_c5\
        );

    \I__883\ : InMux
    port map (
            O => \N__4699\,
            I => \N__4690\
        );

    \I__882\ : InMux
    port map (
            O => \N__4698\,
            I => \N__4690\
        );

    \I__881\ : InMux
    port map (
            O => \N__4697\,
            I => \N__4686\
        );

    \I__880\ : InMux
    port map (
            O => \N__4696\,
            I => \N__4681\
        );

    \I__879\ : InMux
    port map (
            O => \N__4695\,
            I => \N__4681\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__4690\,
            I => \N__4678\
        );

    \I__877\ : InMux
    port map (
            O => \N__4689\,
            I => \N__4675\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__4686\,
            I => \Glue_Lab2_gl_fsm_state_1\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__4681\,
            I => \Glue_Lab2_gl_fsm_state_1\
        );

    \I__874\ : Odrv4
    port map (
            O => \N__4678\,
            I => \Glue_Lab2_gl_fsm_state_1\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__4675\,
            I => \Glue_Lab2_gl_fsm_state_1\
        );

    \I__872\ : InMux
    port map (
            O => \N__4666\,
            I => \N__4663\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__4663\,
            I => \N__4660\
        );

    \I__870\ : Odrv4
    port map (
            O => \N__4660\,
            I => \Glue_Lab2.gl_fsm.enOp_0_a2_2\
        );

    \I__869\ : CascadeMux
    port map (
            O => \N__4657\,
            I => \Glue_Lab2.Gl_subtract_1_cascade_\
        );

    \I__868\ : InMux
    port map (
            O => \N__4654\,
            I => \N__4651\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__4651\,
            I => \N__4648\
        );

    \I__866\ : Odrv12
    port map (
            O => \N__4648\,
            I => \Lab_UT.S_0_s_axbZ0Z3\
        );

    \I__865\ : CascadeMux
    port map (
            O => \N__4645\,
            I => \N__4642\
        );

    \I__864\ : InMux
    port map (
            O => \N__4642\,
            I => \N__4636\
        );

    \I__863\ : InMux
    port map (
            O => \N__4641\,
            I => \N__4636\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__4636\,
            I => \N__4632\
        );

    \I__861\ : InMux
    port map (
            O => \N__4635\,
            I => \N__4629\
        );

    \I__860\ : Odrv4
    port map (
            O => \N__4632\,
            I => \Lab_UT.S_0_s_cZ0Z2\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__4629\,
            I => \Lab_UT.S_0_s_cZ0Z2\
        );

    \I__858\ : CascadeMux
    port map (
            O => \N__4624\,
            I => \Lab_UT.S_m_amZ0Z_2_cascade_\
        );

    \I__857\ : IoInMux
    port map (
            O => \N__4621\,
            I => \N__4618\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__4618\,
            I => \N__4615\
        );

    \I__855\ : Span4Mux_s3_h
    port map (
            O => \N__4615\,
            I => \N__4611\
        );

    \I__854\ : InMux
    port map (
            O => \N__4614\,
            I => \N__4608\
        );

    \I__853\ : Odrv4
    port map (
            O => \N__4611\,
            I => led_c_2
        );

    \I__852\ : LocalMux
    port map (
            O => \N__4608\,
            I => led_c_2
        );

    \I__851\ : InMux
    port map (
            O => \N__4603\,
            I => \N__4598\
        );

    \I__850\ : CascadeMux
    port map (
            O => \N__4602\,
            I => \N__4591\
        );

    \I__849\ : InMux
    port map (
            O => \N__4601\,
            I => \N__4587\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__4598\,
            I => \N__4584\
        );

    \I__847\ : InMux
    port map (
            O => \N__4597\,
            I => \N__4581\
        );

    \I__846\ : InMux
    port map (
            O => \N__4596\,
            I => \N__4578\
        );

    \I__845\ : InMux
    port map (
            O => \N__4595\,
            I => \N__4569\
        );

    \I__844\ : InMux
    port map (
            O => \N__4594\,
            I => \N__4569\
        );

    \I__843\ : InMux
    port map (
            O => \N__4591\,
            I => \N__4569\
        );

    \I__842\ : InMux
    port map (
            O => \N__4590\,
            I => \N__4569\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__4587\,
            I => \Gl_r1_0\
        );

    \I__840\ : Odrv4
    port map (
            O => \N__4584\,
            I => \Gl_r1_0\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__4581\,
            I => \Gl_r1_0\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__4578\,
            I => \Gl_r1_0\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__4569\,
            I => \Gl_r1_0\
        );

    \I__836\ : CascadeMux
    port map (
            O => \N__4558\,
            I => \N__4553\
        );

    \I__835\ : CascadeMux
    port map (
            O => \N__4557\,
            I => \N__4543\
        );

    \I__834\ : InMux
    port map (
            O => \N__4556\,
            I => \N__4532\
        );

    \I__833\ : InMux
    port map (
            O => \N__4553\,
            I => \N__4532\
        );

    \I__832\ : InMux
    port map (
            O => \N__4552\,
            I => \N__4532\
        );

    \I__831\ : InMux
    port map (
            O => \N__4551\,
            I => \N__4532\
        );

    \I__830\ : InMux
    port map (
            O => \N__4550\,
            I => \N__4532\
        );

    \I__829\ : InMux
    port map (
            O => \N__4549\,
            I => \N__4529\
        );

    \I__828\ : InMux
    port map (
            O => \N__4548\,
            I => \N__4523\
        );

    \I__827\ : InMux
    port map (
            O => \N__4547\,
            I => \N__4520\
        );

    \I__826\ : InMux
    port map (
            O => \N__4546\,
            I => \N__4515\
        );

    \I__825\ : InMux
    port map (
            O => \N__4543\,
            I => \N__4515\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__4532\,
            I => \N__4510\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__4529\,
            I => \N__4510\
        );

    \I__822\ : InMux
    port map (
            O => \N__4528\,
            I => \N__4505\
        );

    \I__821\ : InMux
    port map (
            O => \N__4527\,
            I => \N__4505\
        );

    \I__820\ : InMux
    port map (
            O => \N__4526\,
            I => \N__4502\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__4523\,
            I => \Gl_r2_1\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__4520\,
            I => \Gl_r2_1\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__4515\,
            I => \Gl_r2_1\
        );

    \I__816\ : Odrv4
    port map (
            O => \N__4510\,
            I => \Gl_r2_1\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__4505\,
            I => \Gl_r2_1\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__4502\,
            I => \Gl_r2_1\
        );

    \I__813\ : CascadeMux
    port map (
            O => \N__4489\,
            I => \N__4482\
        );

    \I__812\ : CascadeMux
    port map (
            O => \N__4488\,
            I => \N__4479\
        );

    \I__811\ : CascadeMux
    port map (
            O => \N__4487\,
            I => \N__4475\
        );

    \I__810\ : CascadeMux
    port map (
            O => \N__4486\,
            I => \N__4471\
        );

    \I__809\ : InMux
    port map (
            O => \N__4485\,
            I => \N__4468\
        );

    \I__808\ : InMux
    port map (
            O => \N__4482\,
            I => \N__4465\
        );

    \I__807\ : InMux
    port map (
            O => \N__4479\,
            I => \N__4462\
        );

    \I__806\ : InMux
    port map (
            O => \N__4478\,
            I => \N__4453\
        );

    \I__805\ : InMux
    port map (
            O => \N__4475\,
            I => \N__4453\
        );

    \I__804\ : InMux
    port map (
            O => \N__4474\,
            I => \N__4453\
        );

    \I__803\ : InMux
    port map (
            O => \N__4471\,
            I => \N__4453\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__4468\,
            I => \N__4450\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__4465\,
            I => \N__4444\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__4462\,
            I => \N__4444\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__4453\,
            I => \N__4441\
        );

    \I__798\ : Span4Mux_v
    port map (
            O => \N__4450\,
            I => \N__4438\
        );

    \I__797\ : InMux
    port map (
            O => \N__4449\,
            I => \N__4435\
        );

    \I__796\ : Span4Mux_h
    port map (
            O => \N__4444\,
            I => \N__4432\
        );

    \I__795\ : Span4Mux_h
    port map (
            O => \N__4441\,
            I => \N__4429\
        );

    \I__794\ : Odrv4
    port map (
            O => \N__4438\,
            I => \Gl_r2_0\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__4435\,
            I => \Gl_r2_0\
        );

    \I__792\ : Odrv4
    port map (
            O => \N__4432\,
            I => \Gl_r2_0\
        );

    \I__791\ : Odrv4
    port map (
            O => \N__4429\,
            I => \Gl_r2_0\
        );

    \I__790\ : InMux
    port map (
            O => \N__4420\,
            I => \N__4417\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__4417\,
            I => \N__4411\
        );

    \I__788\ : InMux
    port map (
            O => \N__4416\,
            I => \N__4406\
        );

    \I__787\ : InMux
    port map (
            O => \N__4415\,
            I => \N__4406\
        );

    \I__786\ : CascadeMux
    port map (
            O => \N__4414\,
            I => \N__4403\
        );

    \I__785\ : Span4Mux_s2_v
    port map (
            O => \N__4411\,
            I => \N__4391\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__4406\,
            I => \N__4388\
        );

    \I__783\ : InMux
    port map (
            O => \N__4403\,
            I => \N__4385\
        );

    \I__782\ : InMux
    port map (
            O => \N__4402\,
            I => \N__4374\
        );

    \I__781\ : InMux
    port map (
            O => \N__4401\,
            I => \N__4374\
        );

    \I__780\ : InMux
    port map (
            O => \N__4400\,
            I => \N__4374\
        );

    \I__779\ : InMux
    port map (
            O => \N__4399\,
            I => \N__4374\
        );

    \I__778\ : InMux
    port map (
            O => \N__4398\,
            I => \N__4374\
        );

    \I__777\ : InMux
    port map (
            O => \N__4397\,
            I => \N__4367\
        );

    \I__776\ : InMux
    port map (
            O => \N__4396\,
            I => \N__4367\
        );

    \I__775\ : InMux
    port map (
            O => \N__4395\,
            I => \N__4367\
        );

    \I__774\ : InMux
    port map (
            O => \N__4394\,
            I => \N__4364\
        );

    \I__773\ : Odrv4
    port map (
            O => \N__4391\,
            I => \Gl_r1_1\
        );

    \I__772\ : Odrv4
    port map (
            O => \N__4388\,
            I => \Gl_r1_1\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__4385\,
            I => \Gl_r1_1\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__4374\,
            I => \Gl_r1_1\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__4367\,
            I => \Gl_r1_1\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__4364\,
            I => \Gl_r1_1\
        );

    \I__767\ : InMux
    port map (
            O => \N__4351\,
            I => \N__4348\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__4348\,
            I => \Lab_UT.S_m_amZ0Z_1\
        );

    \I__765\ : CascadeMux
    port map (
            O => \N__4345\,
            I => \Lab_UT.S_m_bmZ0Z_1_cascade_\
        );

    \I__764\ : IoInMux
    port map (
            O => \N__4342\,
            I => \N__4339\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__4339\,
            I => \N__4336\
        );

    \I__762\ : Span4Mux_s3_h
    port map (
            O => \N__4336\,
            I => \N__4333\
        );

    \I__761\ : Odrv4
    port map (
            O => \N__4333\,
            I => led_c_1
        );

    \I__760\ : InMux
    port map (
            O => \N__4330\,
            I => \N__4327\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__4327\,
            I => \Glue_Lab2.gl_fsm.enOp_0_a2_1\
        );

    \I__758\ : CascadeMux
    port map (
            O => \N__4324\,
            I => \N__4321\
        );

    \I__757\ : InMux
    port map (
            O => \N__4321\,
            I => \N__4318\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__4318\,
            I => \Glue_Lab2.gl_fsm.enOp_0_a2Z0Z_4\
        );

    \I__755\ : InMux
    port map (
            O => \N__4315\,
            I => \N__4309\
        );

    \I__754\ : InMux
    port map (
            O => \N__4314\,
            I => \N__4304\
        );

    \I__753\ : InMux
    port map (
            O => \N__4313\,
            I => \N__4304\
        );

    \I__752\ : InMux
    port map (
            O => \N__4312\,
            I => \N__4301\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__4309\,
            I => bu_rx_data_rdy
        );

    \I__750\ : LocalMux
    port map (
            O => \N__4304\,
            I => bu_rx_data_rdy
        );

    \I__749\ : LocalMux
    port map (
            O => \N__4301\,
            I => bu_rx_data_rdy
        );

    \I__748\ : CascadeMux
    port map (
            O => \N__4294\,
            I => \Glue_Lab2.Gl_r1_2_1_cascade_\
        );

    \I__747\ : CascadeMux
    port map (
            O => \N__4291\,
            I => \Glue_Lab2.Gl_r1_2_2_cascade_\
        );

    \I__746\ : CascadeMux
    port map (
            O => \N__4288\,
            I => \N__4285\
        );

    \I__745\ : InMux
    port map (
            O => \N__4285\,
            I => \N__4282\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__4282\,
            I => \N__4279\
        );

    \I__743\ : Odrv4
    port map (
            O => \N__4279\,
            I => \Lab_UT.g0Z0Z_1\
        );

    \I__742\ : CascadeMux
    port map (
            O => \N__4276\,
            I => \N__4270\
        );

    \I__741\ : InMux
    port map (
            O => \N__4275\,
            I => \N__4257\
        );

    \I__740\ : InMux
    port map (
            O => \N__4274\,
            I => \N__4257\
        );

    \I__739\ : InMux
    port map (
            O => \N__4273\,
            I => \N__4257\
        );

    \I__738\ : InMux
    port map (
            O => \N__4270\,
            I => \N__4257\
        );

    \I__737\ : InMux
    port map (
            O => \N__4269\,
            I => \N__4257\
        );

    \I__736\ : InMux
    port map (
            O => \N__4268\,
            I => \N__4254\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__4257\,
            I => \Glue_Lab2.enOp\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__4254\,
            I => \Glue_Lab2.enOp\
        );

    \I__733\ : InMux
    port map (
            O => \N__4249\,
            I => \N__4246\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__4246\,
            I => \N__4243\
        );

    \I__731\ : Span4Mux_h
    port map (
            O => \N__4243\,
            I => \N__4240\
        );

    \I__730\ : Odrv4
    port map (
            O => \N__4240\,
            I => \Gl_tx_data_2\
        );

    \I__729\ : InMux
    port map (
            O => \N__4237\,
            I => \N__4234\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__4234\,
            I => \Glue_Lab2.de0.un1_charDataZ0\
        );

    \I__727\ : InMux
    port map (
            O => \N__4231\,
            I => \N__4227\
        );

    \I__726\ : InMux
    port map (
            O => \N__4230\,
            I => \N__4224\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__4227\,
            I => \buart__rx_shifter_fast_5\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__4224\,
            I => \buart__rx_shifter_fast_5\
        );

    \I__723\ : InMux
    port map (
            O => \N__4219\,
            I => \N__4215\
        );

    \I__722\ : InMux
    port map (
            O => \N__4218\,
            I => \N__4212\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__4215\,
            I => \N__4209\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__4212\,
            I => \N__4206\
        );

    \I__719\ : Span4Mux_v
    port map (
            O => \N__4209\,
            I => \N__4201\
        );

    \I__718\ : Span4Mux_s3_h
    port map (
            O => \N__4206\,
            I => \N__4201\
        );

    \I__717\ : Odrv4
    port map (
            O => \N__4201\,
            I => \buart.Z_rx.hhZ0Z_1\
        );

    \I__716\ : InMux
    port map (
            O => \N__4198\,
            I => \N__4195\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__4195\,
            I => \N__4192\
        );

    \I__714\ : Odrv4
    port map (
            O => \N__4192\,
            I => \Glue_Lab2.g0_8_0\
        );

    \I__713\ : InMux
    port map (
            O => \N__4189\,
            I => \N__4186\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__4186\,
            I => \Glue_Lab2.de0.de_escZ0Z_3\
        );

    \I__711\ : CascadeMux
    port map (
            O => \N__4183\,
            I => \N__4174\
        );

    \I__710\ : CascadeMux
    port map (
            O => \N__4182\,
            I => \N__4171\
        );

    \I__709\ : CascadeMux
    port map (
            O => \N__4181\,
            I => \N__4168\
        );

    \I__708\ : CascadeMux
    port map (
            O => \N__4180\,
            I => \N__4165\
        );

    \I__707\ : CascadeMux
    port map (
            O => \N__4179\,
            I => \N__4161\
        );

    \I__706\ : InMux
    port map (
            O => \N__4178\,
            I => \N__4157\
        );

    \I__705\ : InMux
    port map (
            O => \N__4177\,
            I => \N__4154\
        );

    \I__704\ : InMux
    port map (
            O => \N__4174\,
            I => \N__4151\
        );

    \I__703\ : InMux
    port map (
            O => \N__4171\,
            I => \N__4146\
        );

    \I__702\ : InMux
    port map (
            O => \N__4168\,
            I => \N__4146\
        );

    \I__701\ : InMux
    port map (
            O => \N__4165\,
            I => \N__4143\
        );

    \I__700\ : InMux
    port map (
            O => \N__4164\,
            I => \N__4136\
        );

    \I__699\ : InMux
    port map (
            O => \N__4161\,
            I => \N__4136\
        );

    \I__698\ : InMux
    port map (
            O => \N__4160\,
            I => \N__4136\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__4157\,
            I => \buart__rx_bitcount_4\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__4154\,
            I => \buart__rx_bitcount_4\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__4151\,
            I => \buart__rx_bitcount_4\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__4146\,
            I => \buart__rx_bitcount_4\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__4143\,
            I => \buart__rx_bitcount_4\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__4136\,
            I => \buart__rx_bitcount_4\
        );

    \I__691\ : InMux
    port map (
            O => \N__4123\,
            I => \N__4111\
        );

    \I__690\ : InMux
    port map (
            O => \N__4122\,
            I => \N__4108\
        );

    \I__689\ : InMux
    port map (
            O => \N__4121\,
            I => \N__4103\
        );

    \I__688\ : InMux
    port map (
            O => \N__4120\,
            I => \N__4103\
        );

    \I__687\ : InMux
    port map (
            O => \N__4119\,
            I => \N__4096\
        );

    \I__686\ : InMux
    port map (
            O => \N__4118\,
            I => \N__4096\
        );

    \I__685\ : InMux
    port map (
            O => \N__4117\,
            I => \N__4096\
        );

    \I__684\ : InMux
    port map (
            O => \N__4116\,
            I => \N__4089\
        );

    \I__683\ : InMux
    port map (
            O => \N__4115\,
            I => \N__4089\
        );

    \I__682\ : InMux
    port map (
            O => \N__4114\,
            I => \N__4089\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__4111\,
            I => \buart__rx_bitcount_3\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__4108\,
            I => \buart__rx_bitcount_3\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__4103\,
            I => \buart__rx_bitcount_3\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__4096\,
            I => \buart__rx_bitcount_3\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__4089\,
            I => \buart__rx_bitcount_3\
        );

    \I__676\ : CascadeMux
    port map (
            O => \N__4078\,
            I => \buart.Z_rx.bitcount_RNIMK771Z0Z_4_cascade_\
        );

    \I__675\ : InMux
    port map (
            O => \N__4075\,
            I => \N__4069\
        );

    \I__674\ : InMux
    port map (
            O => \N__4074\,
            I => \N__4069\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__4069\,
            I => \buart.Z_rx.idle\
        );

    \I__672\ : CascadeMux
    port map (
            O => \N__4066\,
            I => \buart.Z_rx.idle_cascade_\
        );

    \I__671\ : InMux
    port map (
            O => \N__4063\,
            I => \N__4060\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__4060\,
            I => \N__4056\
        );

    \I__669\ : InMux
    port map (
            O => \N__4059\,
            I => \N__4053\
        );

    \I__668\ : Span4Mux_h
    port map (
            O => \N__4056\,
            I => \N__4050\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__4053\,
            I => \buart.Z_rx.hhZ0Z_0\
        );

    \I__666\ : Odrv4
    port map (
            O => \N__4050\,
            I => \buart.Z_rx.hhZ0Z_0\
        );

    \I__665\ : CascadeMux
    port map (
            O => \N__4045\,
            I => \buart.Z_rx.startbit_cascade_\
        );

    \I__664\ : InMux
    port map (
            O => \N__4042\,
            I => \N__4039\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__4039\,
            I => \buart.Z_rx.bitcount_lm_1\
        );

    \I__662\ : InMux
    port map (
            O => \N__4036\,
            I => \N__4022\
        );

    \I__661\ : InMux
    port map (
            O => \N__4035\,
            I => \N__4022\
        );

    \I__660\ : InMux
    port map (
            O => \N__4034\,
            I => \N__4015\
        );

    \I__659\ : InMux
    port map (
            O => \N__4033\,
            I => \N__4015\
        );

    \I__658\ : InMux
    port map (
            O => \N__4032\,
            I => \N__4015\
        );

    \I__657\ : InMux
    port map (
            O => \N__4031\,
            I => \N__4010\
        );

    \I__656\ : InMux
    port map (
            O => \N__4030\,
            I => \N__4010\
        );

    \I__655\ : InMux
    port map (
            O => \N__4029\,
            I => \N__4003\
        );

    \I__654\ : InMux
    port map (
            O => \N__4028\,
            I => \N__4003\
        );

    \I__653\ : InMux
    port map (
            O => \N__4027\,
            I => \N__4003\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__4022\,
            I => \buart__rx_bitcount_1\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__4015\,
            I => \buart__rx_bitcount_1\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__4010\,
            I => \buart__rx_bitcount_1\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__4003\,
            I => \buart__rx_bitcount_1\
        );

    \I__648\ : InMux
    port map (
            O => \N__3994\,
            I => \N__3991\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__3991\,
            I => \buart.Z_rx.bitcount_cry_1_THRU_CO\
        );

    \I__646\ : InMux
    port map (
            O => \N__3988\,
            I => \N__3980\
        );

    \I__645\ : InMux
    port map (
            O => \N__3987\,
            I => \N__3980\
        );

    \I__644\ : InMux
    port map (
            O => \N__3986\,
            I => \N__3975\
        );

    \I__643\ : InMux
    port map (
            O => \N__3985\,
            I => \N__3975\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__3980\,
            I => \buart.Z_rx.N_29_0_i\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__3975\,
            I => \buart.Z_rx.N_29_0_i\
        );

    \I__640\ : CascadeMux
    port map (
            O => \N__3970\,
            I => \N__3964\
        );

    \I__639\ : InMux
    port map (
            O => \N__3969\,
            I => \N__3957\
        );

    \I__638\ : InMux
    port map (
            O => \N__3968\,
            I => \N__3957\
        );

    \I__637\ : InMux
    port map (
            O => \N__3967\,
            I => \N__3957\
        );

    \I__636\ : InMux
    port map (
            O => \N__3964\,
            I => \N__3954\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__3957\,
            I => \buart.Z_rx.bitcountlde_0\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__3954\,
            I => \buart.Z_rx.bitcountlde_0\
        );

    \I__633\ : CascadeMux
    port map (
            O => \N__3949\,
            I => \buart.Z_rx.bitcount_lm_2_cascade_\
        );

    \I__632\ : InMux
    port map (
            O => \N__3946\,
            I => \N__3937\
        );

    \I__631\ : InMux
    port map (
            O => \N__3945\,
            I => \N__3934\
        );

    \I__630\ : InMux
    port map (
            O => \N__3944\,
            I => \N__3929\
        );

    \I__629\ : InMux
    port map (
            O => \N__3943\,
            I => \N__3929\
        );

    \I__628\ : InMux
    port map (
            O => \N__3942\,
            I => \N__3924\
        );

    \I__627\ : CascadeMux
    port map (
            O => \N__3941\,
            I => \N__3919\
        );

    \I__626\ : CascadeMux
    port map (
            O => \N__3940\,
            I => \N__3916\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__3937\,
            I => \N__3909\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__3934\,
            I => \N__3909\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__3929\,
            I => \N__3909\
        );

    \I__622\ : CascadeMux
    port map (
            O => \N__3928\,
            I => \N__3902\
        );

    \I__621\ : CascadeMux
    port map (
            O => \N__3927\,
            I => \N__3899\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__3924\,
            I => \N__3896\
        );

    \I__619\ : InMux
    port map (
            O => \N__3923\,
            I => \N__3887\
        );

    \I__618\ : InMux
    port map (
            O => \N__3922\,
            I => \N__3887\
        );

    \I__617\ : InMux
    port map (
            O => \N__3919\,
            I => \N__3887\
        );

    \I__616\ : InMux
    port map (
            O => \N__3916\,
            I => \N__3887\
        );

    \I__615\ : Span4Mux_v
    port map (
            O => \N__3909\,
            I => \N__3884\
        );

    \I__614\ : InMux
    port map (
            O => \N__3908\,
            I => \N__3875\
        );

    \I__613\ : InMux
    port map (
            O => \N__3907\,
            I => \N__3875\
        );

    \I__612\ : InMux
    port map (
            O => \N__3906\,
            I => \N__3875\
        );

    \I__611\ : InMux
    port map (
            O => \N__3905\,
            I => \N__3875\
        );

    \I__610\ : InMux
    port map (
            O => \N__3902\,
            I => \N__3872\
        );

    \I__609\ : InMux
    port map (
            O => \N__3899\,
            I => \N__3869\
        );

    \I__608\ : Odrv4
    port map (
            O => \N__3896\,
            I => \buart.Z_rx.startbit\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__3887\,
            I => \buart.Z_rx.startbit\
        );

    \I__606\ : Odrv4
    port map (
            O => \N__3884\,
            I => \buart.Z_rx.startbit\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__3875\,
            I => \buart.Z_rx.startbit\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__3872\,
            I => \buart.Z_rx.startbit\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__3869\,
            I => \buart.Z_rx.startbit\
        );

    \I__602\ : CascadeMux
    port map (
            O => \N__3856\,
            I => \N__3845\
        );

    \I__601\ : CascadeMux
    port map (
            O => \N__3855\,
            I => \N__3841\
        );

    \I__600\ : InMux
    port map (
            O => \N__3854\,
            I => \N__3838\
        );

    \I__599\ : InMux
    port map (
            O => \N__3853\,
            I => \N__3835\
        );

    \I__598\ : InMux
    port map (
            O => \N__3852\,
            I => \N__3832\
        );

    \I__597\ : InMux
    port map (
            O => \N__3851\,
            I => \N__3827\
        );

    \I__596\ : InMux
    port map (
            O => \N__3850\,
            I => \N__3827\
        );

    \I__595\ : InMux
    port map (
            O => \N__3849\,
            I => \N__3822\
        );

    \I__594\ : InMux
    port map (
            O => \N__3848\,
            I => \N__3822\
        );

    \I__593\ : InMux
    port map (
            O => \N__3845\,
            I => \N__3815\
        );

    \I__592\ : InMux
    port map (
            O => \N__3844\,
            I => \N__3815\
        );

    \I__591\ : InMux
    port map (
            O => \N__3841\,
            I => \N__3815\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__3838\,
            I => \buart__rx_bitcount_2\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__3835\,
            I => \buart__rx_bitcount_2\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__3832\,
            I => \buart__rx_bitcount_2\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__3827\,
            I => \buart__rx_bitcount_2\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__3822\,
            I => \buart__rx_bitcount_2\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__3815\,
            I => \buart__rx_bitcount_2\
        );

    \I__584\ : InMux
    port map (
            O => \N__3802\,
            I => \N__3799\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__3799\,
            I => \Glue_Lab2.g0_8_2\
        );

    \I__582\ : InMux
    port map (
            O => \N__3796\,
            I => \N__3793\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__3793\,
            I => \Glue_Lab2.de0.un2_de_hexplusZ0Z_2\
        );

    \I__580\ : CascadeMux
    port map (
            O => \N__3790\,
            I => \Lab_UT.S_0_s_c2_1_cascade_\
        );

    \I__579\ : InMux
    port map (
            O => \N__3787\,
            I => \N__3784\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__3784\,
            I => \Lab_UT.S_0_s_ac0_5_0_2\
        );

    \I__577\ : InMux
    port map (
            O => \N__3781\,
            I => \N__3778\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__3778\,
            I => \N__3775\
        );

    \I__575\ : Odrv4
    port map (
            O => \N__3775\,
            I => \Lab_UT_g1_1\
        );

    \I__574\ : InMux
    port map (
            O => \N__3772\,
            I => \buart.Z_rx.bitcount_cry_0\
        );

    \I__573\ : InMux
    port map (
            O => \N__3769\,
            I => \buart.Z_rx.bitcount_cry_1\
        );

    \I__572\ : InMux
    port map (
            O => \N__3766\,
            I => \buart.Z_rx.bitcount_cry_2\
        );

    \I__571\ : InMux
    port map (
            O => \N__3763\,
            I => \buart.Z_rx.bitcount_cry_3\
        );

    \I__570\ : InMux
    port map (
            O => \N__3760\,
            I => \N__3757\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__3757\,
            I => \buart.Z_rx.bitcount_lm_4\
        );

    \I__568\ : InMux
    port map (
            O => \N__3754\,
            I => \N__3751\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__3751\,
            I => \buart.Z_rx.bitcount_cry_0_THRU_CO\
        );

    \I__566\ : InMux
    port map (
            O => \N__3748\,
            I => \N__3745\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__3745\,
            I => \buart.Z_rx.bitcount_cry_2_THRU_CO\
        );

    \I__564\ : CascadeMux
    port map (
            O => \N__3742\,
            I => \buart.Z_rx.bitcount_lm_3_cascade_\
        );

    \I__563\ : InMux
    port map (
            O => \N__3739\,
            I => \N__3736\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__3736\,
            I => \N__3733\
        );

    \I__561\ : Span4Mux_v
    port map (
            O => \N__3733\,
            I => \N__3730\
        );

    \I__560\ : Odrv4
    port map (
            O => \N__3730\,
            I => \Lab_UT.S_m_bm_N_5LZ0Z7\
        );

    \I__559\ : InMux
    port map (
            O => \N__3727\,
            I => \N__3721\
        );

    \I__558\ : InMux
    port map (
            O => \N__3726\,
            I => \N__3718\
        );

    \I__557\ : InMux
    port map (
            O => \N__3725\,
            I => \N__3713\
        );

    \I__556\ : InMux
    port map (
            O => \N__3724\,
            I => \N__3713\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__3721\,
            I => \Gl_r1_2_rep1\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__3718\,
            I => \Gl_r1_2_rep1\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__3713\,
            I => \Gl_r1_2_rep1\
        );

    \I__552\ : CascadeMux
    port map (
            O => \N__3706\,
            I => \N__3700\
        );

    \I__551\ : CascadeMux
    port map (
            O => \N__3705\,
            I => \N__3697\
        );

    \I__550\ : InMux
    port map (
            O => \N__3704\,
            I => \N__3690\
        );

    \I__549\ : InMux
    port map (
            O => \N__3703\,
            I => \N__3690\
        );

    \I__548\ : InMux
    port map (
            O => \N__3700\,
            I => \N__3690\
        );

    \I__547\ : InMux
    port map (
            O => \N__3697\,
            I => \N__3687\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__3690\,
            I => \N__3684\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__3687\,
            I => \Gl_r2_2_rep1\
        );

    \I__544\ : Odrv4
    port map (
            O => \N__3684\,
            I => \Gl_r2_2_rep1\
        );

    \I__543\ : InMux
    port map (
            O => \N__3679\,
            I => \N__3676\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__3676\,
            I => \Lab_UT.g0_4Z0Z_0\
        );

    \I__541\ : CEMux
    port map (
            O => \N__3673\,
            I => \N__3669\
        );

    \I__540\ : CEMux
    port map (
            O => \N__3672\,
            I => \N__3665\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__3669\,
            I => \N__3662\
        );

    \I__538\ : CEMux
    port map (
            O => \N__3668\,
            I => \N__3659\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__3665\,
            I => \N__3656\
        );

    \I__536\ : Span4Mux_h
    port map (
            O => \N__3662\,
            I => \N__3653\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__3659\,
            I => \N__3650\
        );

    \I__534\ : Span4Mux_v
    port map (
            O => \N__3656\,
            I => \N__3647\
        );

    \I__533\ : Span4Mux_h
    port map (
            O => \N__3653\,
            I => \N__3642\
        );

    \I__532\ : Span4Mux_h
    port map (
            O => \N__3650\,
            I => \N__3642\
        );

    \I__531\ : Odrv4
    port map (
            O => \N__3647\,
            I => \Glue_Lab2.Gl_r17_0_i\
        );

    \I__530\ : Odrv4
    port map (
            O => \N__3642\,
            I => \Glue_Lab2.Gl_r17_0_i\
        );

    \I__529\ : InMux
    port map (
            O => \N__3637\,
            I => \N__3634\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__3634\,
            I => \N__3631\
        );

    \I__527\ : Odrv4
    port map (
            O => \N__3631\,
            I => \Lab_UT.g0_1_0_0\
        );

    \I__526\ : CEMux
    port map (
            O => \N__3628\,
            I => \N__3624\
        );

    \I__525\ : CEMux
    port map (
            O => \N__3627\,
            I => \N__3621\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__3624\,
            I => \Glue_Lab2.Gl_r27_0_i\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__3621\,
            I => \Glue_Lab2.Gl_r27_0_i\
        );

    \I__522\ : InMux
    port map (
            O => \N__3616\,
            I => \N__3613\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__3613\,
            I => \Lab_UT.g0_4_0_0\
        );

    \I__520\ : InMux
    port map (
            O => \N__3610\,
            I => \N__3607\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__3607\,
            I => \Lab_UT.S_1_ac0_1_0Z0Z_0\
        );

    \I__518\ : CascadeMux
    port map (
            O => \N__3604\,
            I => \Lab_UT.S_1_axbZ0Z1_cascade_\
        );

    \I__517\ : InMux
    port map (
            O => \N__3601\,
            I => \N__3598\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__3598\,
            I => \Lab_UT.g1Z0Z_0\
        );

    \I__515\ : CascadeMux
    port map (
            O => \N__3595\,
            I => \Lab_UT.S_0_s_c2_0_cascade_\
        );

    \I__514\ : InMux
    port map (
            O => \N__3592\,
            I => \N__3589\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__3589\,
            I => \Lab_UT.S_0_s_ac0_5_0_1\
        );

    \I__512\ : InMux
    port map (
            O => \N__3586\,
            I => \N__3583\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__3583\,
            I => \Lab_UT.gZ0Z1\
        );

    \I__510\ : CascadeMux
    port map (
            O => \N__3580\,
            I => \N__3576\
        );

    \I__509\ : CascadeMux
    port map (
            O => \N__3579\,
            I => \N__3573\
        );

    \I__508\ : InMux
    port map (
            O => \N__3576\,
            I => \N__3567\
        );

    \I__507\ : InMux
    port map (
            O => \N__3573\,
            I => \N__3567\
        );

    \I__506\ : InMux
    port map (
            O => \N__3572\,
            I => \N__3564\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__3567\,
            I => \Glue_Lab2_Gl_r2_fast_0\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__3564\,
            I => \Glue_Lab2_Gl_r2_fast_0\
        );

    \I__503\ : InMux
    port map (
            O => \N__3559\,
            I => \N__3552\
        );

    \I__502\ : InMux
    port map (
            O => \N__3558\,
            I => \N__3552\
        );

    \I__501\ : CascadeMux
    port map (
            O => \N__3557\,
            I => \N__3549\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__3552\,
            I => \N__3546\
        );

    \I__499\ : InMux
    port map (
            O => \N__3549\,
            I => \N__3543\
        );

    \I__498\ : Odrv4
    port map (
            O => \N__3546\,
            I => \Glue_Lab2_Gl_r1_fast_0\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__3543\,
            I => \Glue_Lab2_Gl_r1_fast_0\
        );

    \I__496\ : CascadeMux
    port map (
            O => \N__3538\,
            I => \Glue_Lab2.gl_fsm.N_14_cascade_\
        );

    \I__495\ : InMux
    port map (
            O => \N__3535\,
            I => \N__3528\
        );

    \I__494\ : InMux
    port map (
            O => \N__3534\,
            I => \N__3528\
        );

    \I__493\ : CascadeMux
    port map (
            O => \N__3533\,
            I => \N__3523\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__3528\,
            I => \N__3519\
        );

    \I__491\ : InMux
    port map (
            O => \N__3527\,
            I => \N__3516\
        );

    \I__490\ : InMux
    port map (
            O => \N__3526\,
            I => \N__3513\
        );

    \I__489\ : InMux
    port map (
            O => \N__3523\,
            I => \N__3508\
        );

    \I__488\ : InMux
    port map (
            O => \N__3522\,
            I => \N__3508\
        );

    \I__487\ : Span4Mux_s2_v
    port map (
            O => \N__3519\,
            I => \N__3503\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__3516\,
            I => \N__3503\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__3513\,
            I => \Glue_Lab2_gl_fsm_state_0\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__3508\,
            I => \Glue_Lab2_gl_fsm_state_0\
        );

    \I__483\ : Odrv4
    port map (
            O => \N__3503\,
            I => \Glue_Lab2_gl_fsm_state_0\
        );

    \I__482\ : InMux
    port map (
            O => \N__3496\,
            I => \N__3493\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__3493\,
            I => \Lab_UT.C_out41_0\
        );

    \I__480\ : CascadeMux
    port map (
            O => \N__3490\,
            I => \led_c_0_4_cascade_\
        );

    \I__479\ : CascadeMux
    port map (
            O => \N__3487\,
            I => \N__3484\
        );

    \I__478\ : InMux
    port map (
            O => \N__3484\,
            I => \N__3481\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__3481\,
            I => \N__3478\
        );

    \I__476\ : Odrv4
    port map (
            O => \N__3478\,
            I => \Gl_tx_data_6\
        );

    \I__475\ : InMux
    port map (
            O => \N__3475\,
            I => \N__3472\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__3472\,
            I => \Lab_UT.S_m_bm_N_2LZ0Z1\
        );

    \I__473\ : IoInMux
    port map (
            O => \N__3469\,
            I => \N__3466\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__3466\,
            I => \N__3463\
        );

    \I__471\ : Span4Mux_s3_h
    port map (
            O => \N__3463\,
            I => \N__3459\
        );

    \I__470\ : InMux
    port map (
            O => \N__3462\,
            I => \N__3456\
        );

    \I__469\ : Odrv4
    port map (
            O => \N__3459\,
            I => led_c_0
        );

    \I__468\ : LocalMux
    port map (
            O => \N__3456\,
            I => led_c_0
        );

    \I__467\ : CascadeMux
    port map (
            O => \N__3451\,
            I => \bu_rx_data_rdy_cascade_\
        );

    \I__466\ : InMux
    port map (
            O => \N__3448\,
            I => \N__3440\
        );

    \I__465\ : InMux
    port map (
            O => \N__3447\,
            I => \N__3437\
        );

    \I__464\ : InMux
    port map (
            O => \N__3446\,
            I => \N__3434\
        );

    \I__463\ : InMux
    port map (
            O => \N__3445\,
            I => \N__3427\
        );

    \I__462\ : InMux
    port map (
            O => \N__3444\,
            I => \N__3427\
        );

    \I__461\ : InMux
    port map (
            O => \N__3443\,
            I => \N__3427\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__3440\,
            I => \N__3424\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__3437\,
            I => \N__3421\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__3434\,
            I => \Glue_Lab2.i_rst_char_detected\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__3427\,
            I => \Glue_Lab2.i_rst_char_detected\
        );

    \I__456\ : Odrv4
    port map (
            O => \N__3424\,
            I => \Glue_Lab2.i_rst_char_detected\
        );

    \I__455\ : Odrv4
    port map (
            O => \N__3421\,
            I => \Glue_Lab2.i_rst_char_detected\
        );

    \I__454\ : CascadeMux
    port map (
            O => \N__3412\,
            I => \N__3409\
        );

    \I__453\ : InMux
    port map (
            O => \N__3409\,
            I => \N__3404\
        );

    \I__452\ : InMux
    port map (
            O => \N__3408\,
            I => \N__3401\
        );

    \I__451\ : InMux
    port map (
            O => \N__3407\,
            I => \N__3398\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__3404\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__3401\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__3398\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__447\ : CascadeMux
    port map (
            O => \N__3391\,
            I => \N__3387\
        );

    \I__446\ : InMux
    port map (
            O => \N__3390\,
            I => \N__3384\
        );

    \I__445\ : InMux
    port map (
            O => \N__3387\,
            I => \N__3381\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__3384\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_5\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__3381\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_5\
        );

    \I__442\ : InMux
    port map (
            O => \N__3376\,
            I => \N__3370\
        );

    \I__441\ : InMux
    port map (
            O => \N__3375\,
            I => \N__3367\
        );

    \I__440\ : InMux
    port map (
            O => \N__3374\,
            I => \N__3362\
        );

    \I__439\ : InMux
    port map (
            O => \N__3373\,
            I => \N__3362\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__3370\,
            I => \N__3359\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__3367\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_3\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__3362\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_3\
        );

    \I__435\ : Odrv4
    port map (
            O => \N__3359\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_3\
        );

    \I__434\ : InMux
    port map (
            O => \N__3352\,
            I => \N__3349\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__3349\,
            I => \N__3346\
        );

    \I__432\ : Odrv4
    port map (
            O => \N__3346\,
            I => \buart.Z_rx.un1_sample_0\
        );

    \I__431\ : CascadeMux
    port map (
            O => \N__3343\,
            I => \buart.Z_rx.ser_clk_2_0_cascade_\
        );

    \I__430\ : CascadeMux
    port map (
            O => \N__3340\,
            I => \Glue_Lab2.de0.un2_de_hexplus_3_xZ0Z0_cascade_\
        );

    \I__429\ : CascadeMux
    port map (
            O => \N__3337\,
            I => \Glue_Lab2.de0.un2_de_hexplus_3_cascade_\
        );

    \I__428\ : CascadeMux
    port map (
            O => \N__3334\,
            I => \Glue_Lab2.is_hexplus_cascade_\
        );

    \I__427\ : InMux
    port map (
            O => \N__3331\,
            I => \N__3328\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__3328\,
            I => \N__3325\
        );

    \I__425\ : Odrv4
    port map (
            O => \N__3325\,
            I => \Gl_tx_data_4\
        );

    \I__424\ : InMux
    port map (
            O => \N__3322\,
            I => \N__3312\
        );

    \I__423\ : InMux
    port map (
            O => \N__3321\,
            I => \N__3312\
        );

    \I__422\ : InMux
    port map (
            O => \N__3320\,
            I => \N__3307\
        );

    \I__421\ : InMux
    port map (
            O => \N__3319\,
            I => \N__3307\
        );

    \I__420\ : InMux
    port map (
            O => \N__3318\,
            I => \N__3304\
        );

    \I__419\ : InMux
    port map (
            O => \N__3317\,
            I => \N__3301\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__3312\,
            I => \buart.Z_rx.ser_clk_2\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__3307\,
            I => \buart.Z_rx.ser_clk_2\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__3304\,
            I => \buart.Z_rx.ser_clk_2\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__3301\,
            I => \buart.Z_rx.ser_clk_2\
        );

    \I__414\ : CascadeMux
    port map (
            O => \N__3292\,
            I => \N__3288\
        );

    \I__413\ : CascadeMux
    port map (
            O => \N__3291\,
            I => \N__3285\
        );

    \I__412\ : InMux
    port map (
            O => \N__3288\,
            I => \N__3280\
        );

    \I__411\ : InMux
    port map (
            O => \N__3285\,
            I => \N__3277\
        );

    \I__410\ : InMux
    port map (
            O => \N__3284\,
            I => \N__3274\
        );

    \I__409\ : InMux
    port map (
            O => \N__3283\,
            I => \N__3271\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__3280\,
            I => \N__3268\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__3277\,
            I => \buart.Z_rx.ser_clk_2_0\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__3274\,
            I => \buart.Z_rx.ser_clk_2_0\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__3271\,
            I => \buart.Z_rx.ser_clk_2_0\
        );

    \I__404\ : Odrv4
    port map (
            O => \N__3268\,
            I => \buart.Z_rx.ser_clk_2_0\
        );

    \I__403\ : CascadeMux
    port map (
            O => \N__3259\,
            I => \N__3255\
        );

    \I__402\ : CascadeMux
    port map (
            O => \N__3258\,
            I => \N__3250\
        );

    \I__401\ : InMux
    port map (
            O => \N__3255\,
            I => \N__3246\
        );

    \I__400\ : InMux
    port map (
            O => \N__3254\,
            I => \N__3241\
        );

    \I__399\ : InMux
    port map (
            O => \N__3253\,
            I => \N__3241\
        );

    \I__398\ : InMux
    port map (
            O => \N__3250\,
            I => \N__3236\
        );

    \I__397\ : InMux
    port map (
            O => \N__3249\,
            I => \N__3236\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__3246\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__3241\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__3236\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__393\ : CascadeMux
    port map (
            O => \N__3229\,
            I => \N__3226\
        );

    \I__392\ : InMux
    port map (
            O => \N__3226\,
            I => \N__3223\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__3223\,
            I => \Glue_Lab2.de0.g0_5_0\
        );

    \I__390\ : InMux
    port map (
            O => \N__3220\,
            I => \N__3217\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__3217\,
            I => \N__3214\
        );

    \I__388\ : Span4Mux_h
    port map (
            O => \N__3214\,
            I => \N__3208\
        );

    \I__387\ : InMux
    port map (
            O => \N__3213\,
            I => \N__3205\
        );

    \I__386\ : InMux
    port map (
            O => \N__3212\,
            I => \N__3200\
        );

    \I__385\ : InMux
    port map (
            O => \N__3211\,
            I => \N__3200\
        );

    \I__384\ : Odrv4
    port map (
            O => \N__3208\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__3205\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__3200\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__381\ : InMux
    port map (
            O => \N__3193\,
            I => \N__3188\
        );

    \I__380\ : InMux
    port map (
            O => \N__3192\,
            I => \N__3185\
        );

    \I__379\ : InMux
    port map (
            O => \N__3191\,
            I => \N__3182\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__3188\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_1\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__3185\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_1\
        );

    \I__376\ : LocalMux
    port map (
            O => \N__3182\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_1\
        );

    \I__375\ : CascadeMux
    port map (
            O => \N__3175\,
            I => \Glue_Lab2.de0.g0_5_2_cascade_\
        );

    \I__374\ : CascadeMux
    port map (
            O => \N__3172\,
            I => \Glue_Lab2.g0_9_2_cascade_\
        );

    \I__373\ : InMux
    port map (
            O => \N__3169\,
            I => \N__3166\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__3166\,
            I => \N__3163\
        );

    \I__371\ : Odrv4
    port map (
            O => \N__3163\,
            I => \Glue_Lab2.g0_7_2\
        );

    \I__370\ : InMux
    port map (
            O => \N__3160\,
            I => \N__3157\
        );

    \I__369\ : LocalMux
    port map (
            O => \N__3157\,
            I => \Glue_Lab2.reset_counte_0_3\
        );

    \I__368\ : CascadeMux
    port map (
            O => \N__3154\,
            I => \buart.Z_rx.bitcount_RNIMK771_0Z0Z_4_cascade_\
        );

    \I__367\ : CascadeMux
    port map (
            O => \N__3151\,
            I => \Glue_Lab2.g0_9_0_cascade_\
        );

    \I__366\ : InMux
    port map (
            O => \N__3148\,
            I => \N__3145\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__3145\,
            I => \Glue_Lab2.reset_counte_0_1\
        );

    \I__364\ : InMux
    port map (
            O => \N__3142\,
            I => \N__3139\
        );

    \I__363\ : LocalMux
    port map (
            O => \N__3139\,
            I => \Glue_Lab2.g0_7_0\
        );

    \I__362\ : CascadeMux
    port map (
            O => \N__3136\,
            I => \buart.Z_rx.bitcountlde_0_cascade_\
        );

    \I__361\ : IoInMux
    port map (
            O => \N__3133\,
            I => \N__3130\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__3130\,
            I => \N__3126\
        );

    \I__359\ : CascadeMux
    port map (
            O => \N__3129\,
            I => \N__3123\
        );

    \I__358\ : Span4Mux_s3_v
    port map (
            O => \N__3126\,
            I => \N__3120\
        );

    \I__357\ : InMux
    port map (
            O => \N__3123\,
            I => \N__3116\
        );

    \I__356\ : Span4Mux_v
    port map (
            O => \N__3120\,
            I => \N__3113\
        );

    \I__355\ : InMux
    port map (
            O => \N__3119\,
            I => \N__3110\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__3116\,
            I => \N__3107\
        );

    \I__353\ : Span4Mux_h
    port map (
            O => \N__3113\,
            I => \N__3104\
        );

    \I__352\ : LocalMux
    port map (
            O => \N__3110\,
            I => \N__3099\
        );

    \I__351\ : Span4Mux_h
    port map (
            O => \N__3107\,
            I => \N__3099\
        );

    \I__350\ : Odrv4
    port map (
            O => \N__3104\,
            I => \CONSTANT_ONE_NET\
        );

    \I__349\ : Odrv4
    port map (
            O => \N__3099\,
            I => \CONSTANT_ONE_NET\
        );

    \I__348\ : CascadeMux
    port map (
            O => \N__3094\,
            I => \buart.Z_rx.N_29_0_i_cascade_\
        );

    \I__347\ : InMux
    port map (
            O => \N__3091\,
            I => \N__3088\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__3088\,
            I => \buart.Z_rx.bitcount_lm_0\
        );

    \I__345\ : CascadeMux
    port map (
            O => \N__3085\,
            I => \N__3082\
        );

    \I__344\ : InMux
    port map (
            O => \N__3082\,
            I => \N__3079\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__3079\,
            I => \N__3076\
        );

    \I__342\ : Odrv12
    port map (
            O => \N__3076\,
            I => \Lab_UT.S_m_bm_N_6LZ0Z10\
        );

    \I__341\ : CascadeMux
    port map (
            O => \N__3073\,
            I => \Lab_UT.g0_0_a3Z0Z_0_cascade_\
        );

    \I__340\ : InMux
    port map (
            O => \N__3070\,
            I => \N__3067\
        );

    \I__339\ : LocalMux
    port map (
            O => \N__3067\,
            I => \Lab_UT.g0_1Z0Z_0\
        );

    \I__338\ : InMux
    port map (
            O => \N__3064\,
            I => \N__3061\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__3061\,
            I => \Lab_UT.N_6\
        );

    \I__336\ : CascadeMux
    port map (
            O => \N__3058\,
            I => \Lab_UT.S_0_s_axbZ0Z3_cascade_\
        );

    \I__335\ : InMux
    port map (
            O => \N__3055\,
            I => \N__3052\
        );

    \I__334\ : LocalMux
    port map (
            O => \N__3052\,
            I => \N__3049\
        );

    \I__333\ : Odrv4
    port map (
            O => \N__3049\,
            I => \Lab_UT.S_m_amZ0Z_3\
        );

    \I__332\ : InMux
    port map (
            O => \N__3046\,
            I => \N__3043\
        );

    \I__331\ : LocalMux
    port map (
            O => \N__3043\,
            I => \N__3040\
        );

    \I__330\ : Odrv12
    port map (
            O => \N__3040\,
            I => \Lab_UT.g1_0_0\
        );

    \I__329\ : CascadeMux
    port map (
            O => \N__3037\,
            I => \Lab_UT.S_m_bmZ0Z_3_cascade_\
        );

    \I__328\ : IoInMux
    port map (
            O => \N__3034\,
            I => \N__3031\
        );

    \I__327\ : LocalMux
    port map (
            O => \N__3031\,
            I => \N__3028\
        );

    \I__326\ : IoSpan4Mux
    port map (
            O => \N__3028\,
            I => \N__3025\
        );

    \I__325\ : Span4Mux_s3_h
    port map (
            O => \N__3025\,
            I => \N__3022\
        );

    \I__324\ : Odrv4
    port map (
            O => \N__3022\,
            I => led_c_3
        );

    \I__323\ : CascadeMux
    port map (
            O => \N__3019\,
            I => \led_c_3_cascade_\
        );

    \I__322\ : InMux
    port map (
            O => \N__3016\,
            I => \N__3013\
        );

    \I__321\ : LocalMux
    port map (
            O => \N__3013\,
            I => \N__3010\
        );

    \I__320\ : Odrv4
    port map (
            O => \N__3010\,
            I => \Gl_tx_data_3\
        );

    \I__319\ : InMux
    port map (
            O => \N__3007\,
            I => \N__3004\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__3004\,
            I => \Lab_UT.S_m_bm_N_3LZ0Z3\
        );

    \I__317\ : CascadeMux
    port map (
            O => \N__3001\,
            I => \Lab_UT.g0_0_a3_0Z0Z_0_cascade_\
        );

    \I__316\ : CascadeMux
    port map (
            O => \N__2998\,
            I => \Lab_UT_C_out41_1_cascade_\
        );

    \I__315\ : InMux
    port map (
            O => \N__2995\,
            I => \N__2992\
        );

    \I__314\ : LocalMux
    port map (
            O => \N__2992\,
            I => \N__2989\
        );

    \I__313\ : Odrv12
    port map (
            O => \N__2989\,
            I => \Gl_tx_data_5\
        );

    \I__312\ : InMux
    port map (
            O => \N__2986\,
            I => \N__2983\
        );

    \I__311\ : LocalMux
    port map (
            O => \N__2983\,
            I => \Lab_UT.N_6_0\
        );

    \I__310\ : InMux
    port map (
            O => \N__2980\,
            I => \N__2977\
        );

    \I__309\ : LocalMux
    port map (
            O => \N__2977\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_ac0_7\
        );

    \I__308\ : CascadeMux
    port map (
            O => \N__2974\,
            I => \buart.Z_rx.ser_clk_2_cascade_\
        );

    \I__307\ : InMux
    port map (
            O => \N__2971\,
            I => \N__2967\
        );

    \I__306\ : InMux
    port map (
            O => \N__2970\,
            I => \N__2964\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__2967\,
            I => \Glue_Lab2.reset_countZ0Z_0\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__2964\,
            I => \Glue_Lab2.reset_countZ0Z_0\
        );

    \I__303\ : InMux
    port map (
            O => \N__2959\,
            I => \N__2956\
        );

    \I__302\ : LocalMux
    port map (
            O => \N__2956\,
            I => \buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_4\
        );

    \I__301\ : InMux
    port map (
            O => \N__2953\,
            I => \N__2950\
        );

    \I__300\ : LocalMux
    port map (
            O => \N__2950\,
            I => \Lab_UT.sDelay.delayRegZ0Z_0\
        );

    \I__299\ : InMux
    port map (
            O => \N__2947\,
            I => \N__2944\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__2944\,
            I => \N__2941\
        );

    \I__297\ : Odrv4
    port map (
            O => \N__2941\,
            I => \Gl_tx_data_0\
        );

    \I__296\ : InMux
    port map (
            O => \N__2938\,
            I => \N__2935\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__2935\,
            I => \buart.Z_tx.shifterZ0Z_2\
        );

    \I__294\ : InMux
    port map (
            O => \N__2932\,
            I => \N__2929\
        );

    \I__293\ : LocalMux
    port map (
            O => \N__2929\,
            I => \buart.Z_tx.shifterZ0Z_3\
        );

    \I__292\ : InMux
    port map (
            O => \N__2926\,
            I => \N__2923\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__2923\,
            I => \buart.Z_tx.shifterZ0Z_4\
        );

    \I__290\ : InMux
    port map (
            O => \N__2920\,
            I => \N__2917\
        );

    \I__289\ : LocalMux
    port map (
            O => \N__2917\,
            I => \buart.Z_tx.shifterZ0Z_5\
        );

    \I__288\ : InMux
    port map (
            O => \N__2914\,
            I => \N__2911\
        );

    \I__287\ : LocalMux
    port map (
            O => \N__2911\,
            I => \buart.Z_tx.shifterZ0Z_7\
        );

    \I__286\ : InMux
    port map (
            O => \N__2908\,
            I => \N__2905\
        );

    \I__285\ : LocalMux
    port map (
            O => \N__2905\,
            I => \buart.Z_tx.shifterZ0Z_6\
        );

    \I__284\ : InMux
    port map (
            O => \N__2902\,
            I => \N__2899\
        );

    \I__283\ : LocalMux
    port map (
            O => \N__2899\,
            I => \Glue_Lab2.reset_count_cry_2_THRU_CO\
        );

    \I__282\ : CascadeMux
    port map (
            O => \N__2896\,
            I => \N__2893\
        );

    \I__281\ : InMux
    port map (
            O => \N__2893\,
            I => \N__2889\
        );

    \I__280\ : InMux
    port map (
            O => \N__2892\,
            I => \N__2886\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__2889\,
            I => \Glue_Lab2.reset_countZ0Z_3\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__2886\,
            I => \Glue_Lab2.reset_countZ0Z_3\
        );

    \I__277\ : CascadeMux
    port map (
            O => \N__2881\,
            I => \N__2878\
        );

    \I__276\ : InMux
    port map (
            O => \N__2878\,
            I => \N__2875\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__2875\,
            I => \Glue_Lab2.reset_count_cry_0_THRU_CO\
        );

    \I__274\ : InMux
    port map (
            O => \N__2872\,
            I => \N__2868\
        );

    \I__273\ : InMux
    port map (
            O => \N__2871\,
            I => \N__2865\
        );

    \I__272\ : LocalMux
    port map (
            O => \N__2868\,
            I => \Glue_Lab2.reset_countZ0Z_1\
        );

    \I__271\ : LocalMux
    port map (
            O => \N__2865\,
            I => \Glue_Lab2.reset_countZ0Z_1\
        );

    \I__270\ : CascadeMux
    port map (
            O => \N__2860\,
            I => \buart.Z_rx.Z_baudgen.counter_0_1_5_cascade_\
        );

    \I__269\ : InMux
    port map (
            O => \N__2857\,
            I => \Glue_Lab2.reset_count_cry_1\
        );

    \I__268\ : InMux
    port map (
            O => \N__2854\,
            I => \Glue_Lab2.reset_count_cry_2\
        );

    \I__267\ : InMux
    port map (
            O => \N__2851\,
            I => \Glue_Lab2.reset_count_cry_3\
        );

    \I__266\ : InMux
    port map (
            O => \N__2848\,
            I => \N__2845\
        );

    \I__265\ : LocalMux
    port map (
            O => \N__2845\,
            I => \N__2842\
        );

    \I__264\ : Odrv4
    port map (
            O => \N__2842\,
            I => \Glue_Lab2.reset_count_cry_1_THRU_CO\
        );

    \I__263\ : CascadeMux
    port map (
            O => \N__2839\,
            I => \N__2835\
        );

    \I__262\ : CascadeMux
    port map (
            O => \N__2838\,
            I => \N__2832\
        );

    \I__261\ : InMux
    port map (
            O => \N__2835\,
            I => \N__2829\
        );

    \I__260\ : InMux
    port map (
            O => \N__2832\,
            I => \N__2826\
        );

    \I__259\ : LocalMux
    port map (
            O => \N__2829\,
            I => \N__2823\
        );

    \I__258\ : LocalMux
    port map (
            O => \N__2826\,
            I => \Glue_Lab2.reset_countZ0Z_2\
        );

    \I__257\ : Odrv4
    port map (
            O => \N__2823\,
            I => \Glue_Lab2.reset_countZ0Z_2\
        );

    \I__256\ : InMux
    port map (
            O => \N__2818\,
            I => \N__2815\
        );

    \I__255\ : LocalMux
    port map (
            O => \N__2815\,
            I => \buart.Z_tx.shifterZ0Z_1\
        );

    \I__254\ : InMux
    port map (
            O => \N__2812\,
            I => \N__2809\
        );

    \I__253\ : LocalMux
    port map (
            O => \N__2809\,
            I => \buart.Z_tx.shifterZ0Z_0\
        );

    \I__252\ : IoInMux
    port map (
            O => \N__2806\,
            I => \N__2803\
        );

    \I__251\ : LocalMux
    port map (
            O => \N__2803\,
            I => \N__2800\
        );

    \I__250\ : IoSpan4Mux
    port map (
            O => \N__2800\,
            I => \N__2797\
        );

    \I__249\ : Odrv4
    port map (
            O => \N__2797\,
            I => clk_in_c
        );

    \I__248\ : IoInMux
    port map (
            O => \N__2794\,
            I => \N__2791\
        );

    \I__247\ : LocalMux
    port map (
            O => \N__2791\,
            I => \N__2788\
        );

    \I__246\ : Span4Mux_s1_h
    port map (
            O => \N__2788\,
            I => \N__2785\
        );

    \I__245\ : Span4Mux_h
    port map (
            O => \N__2785\,
            I => \N__2782\
        );

    \I__244\ : Sp12to4
    port map (
            O => \N__2782\,
            I => \N__2779\
        );

    \I__243\ : Odrv12
    port map (
            O => \N__2779\,
            I => clk
        );

    \I__242\ : InMux
    port map (
            O => \N__2776\,
            I => \N__2773\
        );

    \I__241\ : LocalMux
    port map (
            O => \N__2773\,
            I => \N__2770\
        );

    \I__240\ : Span4Mux_h
    port map (
            O => \N__2770\,
            I => \N__2767\
        );

    \I__239\ : IoSpan4Mux
    port map (
            O => \N__2767\,
            I => \N__2764\
        );

    \I__238\ : Odrv4
    port map (
            O => \N__2764\,
            I => \uart_RXD\
        );

    \I__237\ : IoInMux
    port map (
            O => \N__2761\,
            I => \N__2758\
        );

    \I__236\ : LocalMux
    port map (
            O => \N__2758\,
            I => \N__2755\
        );

    \I__235\ : IoSpan4Mux
    port map (
            O => \N__2755\,
            I => \N__2752\
        );

    \I__234\ : Span4Mux_s3_h
    port map (
            O => \N__2752\,
            I => \N__2749\
        );

    \I__233\ : Odrv4
    port map (
            O => \N__2749\,
            I => o_serial_data_c
        );

    \I__232\ : InMux
    port map (
            O => \N__2746\,
            I => \Glue_Lab2.reset_count_cry_0\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_9_0_\
        );

    \IN_MUX_bfv_6_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_11_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \clk_derived_clock_RNI7BQ7\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2794\,
            GLOBALBUFFEROUTPUT => clk_g
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \buart.Z_rx.hh_1_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4059\,
            lcout => \buart.Z_rx.hhZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6163\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.hh_0_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2776\,
            lcout => \buart.Z_rx.hhZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6163\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.uart_tx_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2812\,
            in2 => \_gnd_net_\,
            in3 => \N__6796\,
            lcout => o_serial_data_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6165\,
            ce => \N__6711\,
            sr => \_gnd_net_\
        );

    \Glue_Lab2.reset_count_cry_c_0_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2970\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_11_0_\,
            carryout => \Glue_Lab2.reset_count_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.reset_count_cry_0_THRU_LUT4_0_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2871\,
            in2 => \_gnd_net_\,
            in3 => \N__2746\,
            lcout => \Glue_Lab2.reset_count_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \Glue_Lab2.reset_count_cry_0\,
            carryout => \Glue_Lab2.reset_count_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.reset_count_cry_1_THRU_LUT4_0_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2839\,
            in3 => \N__2857\,
            lcout => \Glue_Lab2.reset_count_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \Glue_Lab2.reset_count_cry_1\,
            carryout => \Glue_Lab2.reset_count_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.reset_count_cry_2_THRU_LUT4_0_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2892\,
            in2 => \_gnd_net_\,
            in3 => \N__2854\,
            lcout => \Glue_Lab2.reset_count_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \Glue_Lab2.reset_count_cry_2\,
            carryout => \Glue_Lab2.reset_count_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.reset_count_4_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__3447\,
            in1 => \N__5292\,
            in2 => \_gnd_net_\,
            in3 => \N__2851\,
            lcout => \Glue_Lab2.reset_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6166\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_0_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3213\,
            in2 => \_gnd_net_\,
            in3 => \N__3946\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6166\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.reset_count_2_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011010010"
        )
    port map (
            in0 => \N__2848\,
            in1 => \N__3148\,
            in2 => \N__2838\,
            in3 => \N__3448\,
            lcout => \Glue_Lab2.reset_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6164\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_1_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__6789\,
            in1 => \N__2938\,
            in2 => \_gnd_net_\,
            in3 => \N__2947\,
            lcout => \buart.Z_tx.shifterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6167\,
            ce => \N__6715\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_0_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6788\,
            in2 => \_gnd_net_\,
            in3 => \N__2818\,
            lcout => \buart.Z_tx.shifterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6167\,
            ce => \N__6715\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_7_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__6795\,
            in1 => \_gnd_net_\,
            in2 => \N__3487\,
            in3 => \N__6727\,
            lcout => \buart.Z_tx.shifterZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6167\,
            ce => \N__6715\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_2_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__2932\,
            in1 => \N__6790\,
            in2 => \_gnd_net_\,
            in3 => \N__4762\,
            lcout => \buart.Z_tx.shifterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6167\,
            ce => \N__6715\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_3_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__6791\,
            in1 => \N__2926\,
            in2 => \_gnd_net_\,
            in3 => \N__4249\,
            lcout => \buart.Z_tx.shifterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6167\,
            ce => \N__6715\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_4_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__2920\,
            in1 => \N__6792\,
            in2 => \_gnd_net_\,
            in3 => \N__3016\,
            lcout => \buart.Z_tx.shifterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6167\,
            ce => \N__6715\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_5_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6793\,
            in1 => \N__3331\,
            in2 => \_gnd_net_\,
            in3 => \N__2908\,
            lcout => \buart.Z_tx.shifterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6167\,
            ce => \N__6715\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_6_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__2914\,
            in1 => \N__6794\,
            in2 => \_gnd_net_\,
            in3 => \N__2995\,
            lcout => \buart.Z_tx.shifterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6167\,
            ce => \N__6715\,
            sr => \_gnd_net_\
        );

    \Glue_Lab2.reset_count_3_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000010100"
        )
    port map (
            in0 => \N__3443\,
            in1 => \N__2902\,
            in2 => \N__2896\,
            in3 => \N__5248\,
            lcout => \Glue_Lab2.reset_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6168\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.reset_count_1_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010011010"
        )
    port map (
            in0 => \N__2872\,
            in1 => \N__5509\,
            in2 => \N__2881\,
            in3 => \N__3445\,
            lcout => \Glue_Lab2.reset_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6168\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNO_0_5_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__3212\,
            in1 => \N__3192\,
            in2 => \_gnd_net_\,
            in3 => \N__3283\,
            lcout => OPEN,
            ltout => \buart.Z_rx.Z_baudgen.counter_0_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_5_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100000"
        )
    port map (
            in0 => \N__3390\,
            in1 => \N__2980\,
            in2 => \N__2860\,
            in3 => \N__3945\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6168\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNO_1_5_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3374\,
            in1 => \N__3254\,
            in2 => \N__3412\,
            in3 => \N__3318\,
            lcout => \buart.Z_rx.Z_baudgen.un5_counter_ac0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNIT3N1_1_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3191\,
            in2 => \_gnd_net_\,
            in3 => \N__3211\,
            lcout => \buart.Z_rx.ser_clk_2\,
            ltout => \buart.Z_rx.ser_clk_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNO_0_4_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__3373\,
            in1 => \N__3408\,
            in2 => \N__2974\,
            in3 => \N__3253\,
            lcout => \buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.reset_count_0_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010011010"
        )
    port map (
            in0 => \N__2971\,
            in1 => \N__3160\,
            in2 => \N__3129\,
            in3 => \N__3444\,
            lcout => \Glue_Lab2.reset_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6168\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.sDelay.delayReg_1_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__2953\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6247\,
            lcout => \Lab_UT.sDelay.delayRegZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_4_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010001000100"
        )
    port map (
            in0 => \N__3943\,
            in1 => \N__2959\,
            in2 => \N__3291\,
            in3 => \N__3321\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_3_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__3322\,
            in1 => \N__3375\,
            in2 => \N__3259\,
            in3 => \N__3944\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.sDelay.delayReg_0_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6246\,
            in1 => \N__4697\,
            in2 => \_gnd_net_\,
            in3 => \N__3526\,
            lcout => \Lab_UT.sDelay.delayRegZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_tx_data_0_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__3462\,
            in1 => \N__5382\,
            in2 => \_gnd_net_\,
            in3 => \N__5016\,
            lcout => \Gl_tx_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_rst_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__5293\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3446\,
            lcout => \Gl_rst\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.S_m_bm_3_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001100011"
        )
    port map (
            in0 => \N__3739\,
            in1 => \N__3007\,
            in2 => \N__3085\,
            in3 => \N__3475\,
            lcout => OPEN,
            ltout => \Lab_UT.S_m_bmZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.S_m_ns_3_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3055\,
            in2 => \N__3037\,
            in3 => \N__5571\,
            lcout => led_c_3,
            ltout => \led_c_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_tx_data_3_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6614\,
            in2 => \N__3019\,
            in3 => \N__5017\,
            lcout => \Gl_tx_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6173\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.S_m_bm_N_3L3_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5651\,
            in2 => \_gnd_net_\,
            in3 => \N__5718\,
            lcout => \Lab_UT.S_m_bm_N_3LZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.g0_0_a3_0_1_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100100011"
        )
    port map (
            in0 => \N__5720\,
            in1 => \N__5813\,
            in2 => \N__5661\,
            in3 => \N__5882\,
            lcout => OPEN,
            ltout => \Lab_UT.g0_0_a3_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.g0_1_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__3637\,
            in1 => \N__3046\,
            in2 => \N__3001\,
            in3 => \N__2986\,
            lcout => OPEN,
            ltout => \Lab_UT_C_out41_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_tx_data_5_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111010001"
        )
    port map (
            in0 => \N__3781\,
            in1 => \N__5896\,
            in2 => \N__2998\,
            in3 => \N__5018\,
            lcout => \Gl_tx_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6173\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.g0_0_a3_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5652\,
            in2 => \_gnd_net_\,
            in3 => \N__5719\,
            lcout => \Lab_UT.N_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_r1_1_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__6352\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6474\,
            lcout => \Gl_r1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6178\,
            ce => \N__3668\,
            sr => \_gnd_net_\
        );

    \Lab_UT.g0_0_a3_0_0_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100100011"
        )
    port map (
            in0 => \N__5717\,
            in1 => \N__3704\,
            in2 => \N__5656\,
            in3 => \N__3725\,
            lcout => OPEN,
            ltout => \Lab_UT.g0_0_a3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.g0_0_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__3601\,
            in1 => \N__3070\,
            in2 => \N__3073\,
            in3 => \N__3064\,
            lcout => \Lab_UT.C_out41_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.g0_1_0_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111010"
        )
    port map (
            in0 => \N__3726\,
            in1 => \N__4549\,
            in2 => \N__4414\,
            in3 => \N__3703\,
            lcout => \Lab_UT.g0_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.g0_0_a3_0_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5642\,
            in2 => \_gnd_net_\,
            in3 => \N__5715\,
            lcout => \Lab_UT.N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_r1_3_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6353\,
            in2 => \_gnd_net_\,
            in3 => \N__6615\,
            lcout => \Gl_r1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6178\,
            ce => \N__3668\,
            sr => \_gnd_net_\
        );

    \Lab_UT.g0_3_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010000000"
        )
    port map (
            in0 => \N__3724\,
            in1 => \N__5641\,
            in2 => \N__3706\,
            in3 => \N__5716\,
            lcout => \Lab_UT.S_0_s_ac0_5_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.S_0_s_axb3_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5633\,
            in2 => \_gnd_net_\,
            in3 => \N__5721\,
            lcout => \Lab_UT.S_0_s_axbZ0Z3\,
            ltout => \Lab_UT.S_0_s_axbZ0Z3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.S_m_am_3_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111001111000"
        )
    port map (
            in0 => \N__5784\,
            in1 => \N__5863\,
            in2 => \N__3058\,
            in3 => \N__4635\,
            lcout => \Lab_UT.S_m_amZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.g1_2_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101001000101"
        )
    port map (
            in0 => \N__4397\,
            in1 => \N__4596\,
            in2 => \N__4489\,
            in3 => \N__4547\,
            lcout => \Lab_UT.g1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.gl_fsm.state_RNITO9T5_0_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__3535\,
            in1 => \N__4699\,
            in2 => \N__6361\,
            in3 => \N__5031\,
            lcout => \Glue_Lab2.Gl_r27_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.g0_4_1_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001001001000"
        )
    port map (
            in0 => \N__5864\,
            in1 => \N__5632\,
            in2 => \N__5811\,
            in3 => \N__5722\,
            lcout => \Lab_UT.g0_4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.S_m_bm_N_6L10_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__3559\,
            in1 => \N__4528\,
            in2 => \N__3580\,
            in3 => \N__4396\,
            lcout => \Lab_UT.S_m_bm_N_6LZ0Z10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.gl_fsm.state_RNITO9T5_0_0_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__4698\,
            in1 => \N__6348\,
            in2 => \N__5037\,
            in3 => \N__3534\,
            lcout => \Glue_Lab2.Gl_r17_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.S_0_s_c2_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010000000"
        )
    port map (
            in0 => \N__3558\,
            in1 => \N__4527\,
            in2 => \N__3579\,
            in3 => \N__4395\,
            lcout => \Lab_UT.S_0_s_cZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_r2_fast_0_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5388\,
            in2 => \_gnd_net_\,
            in3 => \N__6358\,
            lcout => \Glue_Lab2_Gl_r2_fast_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6188\,
            ce => \N__3627\,
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_r2_fast_2_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5227\,
            in2 => \_gnd_net_\,
            in3 => \N__6357\,
            lcout => \Gl_r2_fast_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6188\,
            ce => \N__3627\,
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_r2_2_rep1_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__6355\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5228\,
            lcout => \Gl_r2_2_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6188\,
            ce => \N__3627\,
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_r2_3_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6356\,
            in2 => \_gnd_net_\,
            in3 => \N__6619\,
            lcout => \Gl_r2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6188\,
            ce => \N__3627\,
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_r2_0_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__5389\,
            in1 => \N__6354\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Gl_r2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6188\,
            ce => \N__3627\,
            sr => \_gnd_net_\
        );

    \Glue_Lab2.de0.g0_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__5229\,
            in1 => \N__5439\,
            in2 => \N__3229\,
            in3 => \N__5387\,
            lcout => OPEN,
            ltout => \Glue_Lab2.g0_9_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.reset_count_RNO_0_2_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__4198\,
            in1 => \N__5305\,
            in2 => \N__3151\,
            in3 => \N__3142\,
            lcout => \Glue_Lab2.reset_counte_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.de0.g0_4_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__4117\,
            in1 => \N__3848\,
            in2 => \N__4181\,
            in3 => \N__4032\,
            lcout => \Glue_Lab2.g0_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.de0.g0_0_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__4119\,
            in1 => \N__3849\,
            in2 => \N__4182\,
            in3 => \N__4034\,
            lcout => \Glue_Lab2.g0_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.de0.g0_12_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__4033\,
            in1 => \N__4118\,
            in2 => \N__4183\,
            in3 => \N__3852\,
            lcout => \Glue_Lab2.g0_7_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_4_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100100000"
        )
    port map (
            in0 => \N__4178\,
            in1 => \N__3907\,
            in2 => \N__3970\,
            in3 => \N__3760\,
            lcout => \buart__rx_bitcount_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6169\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNILM873_0_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011111"
        )
    port map (
            in0 => \N__3317\,
            in1 => \N__4075\,
            in2 => \N__3292\,
            in3 => \N__4314\,
            lcout => \buart.Z_rx.bitcountlde_0\,
            ltout => \buart.Z_rx.bitcountlde_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_0_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100100000"
        )
    port map (
            in0 => \N__5447\,
            in1 => \N__3906\,
            in2 => \N__3136\,
            in3 => \N__3091\,
            lcout => \buart__rx_bitcount_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6169\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNIIU223_0_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4313\,
            in2 => \_gnd_net_\,
            in3 => \N__4074\,
            lcout => \buart.Z_rx.N_29_0_i\,
            ltout => \buart.Z_rx.N_29_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNO_0_0_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011011110110"
        )
    port map (
            in0 => \N__3119\,
            in1 => \N__5443\,
            in2 => \N__3094\,
            in3 => \N__3905\,
            lcout => \buart.Z_rx.bitcount_lm_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.de0.g0_2_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__5099\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6091\,
            lcout => \Glue_Lab2.de0.g0_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_1_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__3193\,
            in1 => \N__3220\,
            in2 => \_gnd_net_\,
            in3 => \N__3908\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6169\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNIMK771_1_4_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4028\,
            in1 => \N__4115\,
            in2 => \N__4179\,
            in3 => \N__3844\,
            lcout => \buart.Z_rx.un1_sample_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.de0.g0_7_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__4116\,
            in1 => \N__4164\,
            in2 => \N__3856\,
            in3 => \N__4029\,
            lcout => \Glue_Lab2.g0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.de0.g0_14_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5104\,
            in2 => \_gnd_net_\,
            in3 => \N__5499\,
            lcout => OPEN,
            ltout => \Glue_Lab2.de0.g0_5_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.de0.g0_11_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__5436\,
            in1 => \N__5230\,
            in2 => \N__3175\,
            in3 => \N__5355\,
            lcout => OPEN,
            ltout => \Glue_Lab2.g0_9_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.reset_count_RNO_0_0_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__5294\,
            in1 => \N__3802\,
            in2 => \N__3172\,
            in3 => \N__3169\,
            lcout => \Glue_Lab2.reset_counte_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNIMK771_0_4_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__4114\,
            in1 => \N__4027\,
            in2 => \N__3855\,
            in3 => \N__4160\,
            lcout => OPEN,
            ltout => \buart.Z_rx.bitcount_RNIMK771_0Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNI9F1H1_0_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3154\,
            in3 => \N__5435\,
            lcout => bu_rx_data_rdy,
            ltout => \bu_rx_data_rdy_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.de0.de_esc_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4900\,
            in1 => \N__4189\,
            in2 => \N__3451\,
            in3 => \N__5356\,
            lcout => \Glue_Lab2.i_rst_char_detected\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNI6KE3_5_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__3249\,
            in1 => \N__3407\,
            in2 => \N__3391\,
            in3 => \N__3376\,
            lcout => \buart.Z_rx.ser_clk_2_0\,
            ltout => \buart.Z_rx.ser_clk_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNIC77M1_0_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__3352\,
            in1 => \N__3319\,
            in2 => \N__3343\,
            in3 => \N__5453\,
            lcout => \buart.Z_rx.sample\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.de0.un2_de_hexplus_3_x0_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__4231\,
            in1 => \N__5196\,
            in2 => \N__6471\,
            in3 => \N__5344\,
            lcout => OPEN,
            ltout => \Glue_Lab2.de0.un2_de_hexplus_3_xZ0Z0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.de0.un2_de_hexplus_3_ns_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3340\,
            in3 => \N__6090\,
            lcout => OPEN,
            ltout => \Glue_Lab2.de0.un2_de_hexplus_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.de0.de_hexplus_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__3796\,
            in1 => \N__4237\,
            in2 => \N__3337\,
            in3 => \N__4312\,
            lcout => \Glue_Lab2.is_hexplus\,
            ltout => \Glue_Lab2.is_hexplus_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_tx_data_4_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110101111"
        )
    port map (
            in0 => \N__5500\,
            in1 => \_gnd_net_\,
            in2 => \N__3334\,
            in3 => \_gnd_net_\,
            lcout => \Gl_tx_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6174\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_2_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010010"
        )
    port map (
            in0 => \N__3320\,
            in1 => \N__3284\,
            in2 => \N__3258\,
            in3 => \N__3942\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6174\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.gl_fsm.state_RNIDFRT_0_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000100000"
        )
    port map (
            in0 => \N__5345\,
            in1 => \N__3527\,
            in2 => \N__6469\,
            in3 => \N__5197\,
            lcout => \Glue_Lab2.gl_fsm.enOp_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.gl_fsm.state_1_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100100000"
        )
    port map (
            in0 => \N__5010\,
            in1 => \N__6249\,
            in2 => \N__3533\,
            in3 => \N__4696\,
            lcout => \Glue_Lab2_gl_fsm_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6179\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.gl_fsm.state_ns_1_0__m1_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3522\,
            in2 => \_gnd_net_\,
            in3 => \N__5008\,
            lcout => OPEN,
            ltout => \Glue_Lab2.gl_fsm.N_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.gl_fsm.state_0_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__6248\,
            in1 => \N__4695\,
            in2 => \N__3538\,
            in3 => \N__4268\,
            lcout => \Glue_Lab2_gl_fsm_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6179\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.g0_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110011101100"
        )
    port map (
            in0 => \N__5950\,
            in1 => \N__3586\,
            in2 => \N__4288\,
            in3 => \N__3496\,
            lcout => OPEN,
            ltout => \led_c_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_tx_data_6_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__5009\,
            in1 => \_gnd_net_\,
            in2 => \N__3490\,
            in3 => \N__5130\,
            lcout => \Gl_tx_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6179\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.S_m_bm_N_2L1_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5800\,
            in2 => \_gnd_net_\,
            in3 => \N__5873\,
            lcout => \Lab_UT.S_m_bm_N_2LZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.S_m_0_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__4601\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4485\,
            lcout => led_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.S_1_ac0_1_0_0_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001100"
        )
    port map (
            in0 => \N__5805\,
            in1 => \N__4401\,
            in2 => \N__4558\,
            in3 => \N__5872\,
            lcout => \Lab_UT.S_1_ac0_1_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.S_1_axb1_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__4402\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4556\,
            lcout => OPEN,
            ltout => \Lab_UT.S_1_axbZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.S_1_ac0_1_0_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011111100"
        )
    port map (
            in0 => \N__4595\,
            in1 => \N__3610\,
            in2 => \N__3604\,
            in3 => \N__4478\,
            lcout => \Lab_UT.S_1_c3_d\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.S_m_am_1_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010101101010"
        )
    port map (
            in0 => \N__4400\,
            in1 => \N__4594\,
            in2 => \N__4487\,
            in3 => \N__4552\,
            lcout => \Lab_UT.S_m_amZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_r1_0_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6291\,
            in2 => \_gnd_net_\,
            in3 => \N__5383\,
            lcout => \Gl_r1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6185\,
            ce => \N__3673\,
            sr => \_gnd_net_\
        );

    \Lab_UT.g1_0_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101001000101"
        )
    port map (
            in0 => \N__4398\,
            in1 => \N__4590\,
            in2 => \N__4486\,
            in3 => \N__4550\,
            lcout => \Lab_UT.g1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.g0_7_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100010001000"
        )
    port map (
            in0 => \N__4551\,
            in1 => \N__4399\,
            in2 => \N__4602\,
            in3 => \N__4474\,
            lcout => OPEN,
            ltout => \Lab_UT.S_0_s_c2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.g1_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3679\,
            in2 => \N__3595\,
            in3 => \N__3592\,
            lcout => \Lab_UT.gZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.S_m_bm_1_2_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110101000100"
        )
    port map (
            in0 => \N__4394\,
            in1 => \N__4526\,
            in2 => \N__3557\,
            in3 => \N__3572\,
            lcout => \Lab_UT.S_m_bm_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_r1_fast_0_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6359\,
            in3 => \N__5386\,
            lcout => \Glue_Lab2_Gl_r1_fast_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6189\,
            ce => \N__3672\,
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_r1_fast_2_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__5234\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6343\,
            lcout => \Gl_r1_fast_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6189\,
            ce => \N__3672\,
            sr => \_gnd_net_\
        );

    \Lab_UT.S_m_bm_N_5L7_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__4746\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4734\,
            lcout => \Lab_UT.S_m_bm_N_5LZ0Z7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_r1_2_rep1_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__5233\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6339\,
            lcout => \Gl_r1_2_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6189\,
            ce => \N__3672\,
            sr => \_gnd_net_\
        );

    \Lab_UT.g0_4_0_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001001001000"
        )
    port map (
            in0 => \N__3727\,
            in1 => \N__5631\,
            in2 => \N__3705\,
            in3 => \N__5723\,
            lcout => \Lab_UT.g0_4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_r1_2_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__5232\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6338\,
            lcout => \Gl_r1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6189\,
            ce => \N__3672\,
            sr => \_gnd_net_\
        );

    \Lab_UT.g0_4_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010000000"
        )
    port map (
            in0 => \N__5860\,
            in1 => \N__5630\,
            in2 => \N__5801\,
            in3 => \N__5724\,
            lcout => \Lab_UT.S_0_s_ac0_5_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.g0_1_1_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100001010"
        )
    port map (
            in0 => \N__5871\,
            in1 => \N__4546\,
            in2 => \N__5812\,
            in3 => \N__4416\,
            lcout => \Lab_UT.g0_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_r2_1_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6344\,
            in2 => \_gnd_net_\,
            in3 => \N__6475\,
            lcout => \Gl_r2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6192\,
            ce => \N__3628\,
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_r2_2_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__5235\,
            in1 => \_gnd_net_\,
            in2 => \N__6360\,
            in3 => \_gnd_net_\,
            lcout => \Gl_r2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6192\,
            ce => \N__3628\,
            sr => \_gnd_net_\
        );

    \Lab_UT.g0_2_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100010100000"
        )
    port map (
            in0 => \N__4415\,
            in1 => \N__4449\,
            in2 => \N__4557\,
            in3 => \N__4603\,
            lcout => OPEN,
            ltout => \Lab_UT.S_0_s_c2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.g1_1_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3616\,
            in2 => \N__3790\,
            in3 => \N__3787\,
            lcout => \Lab_UT_g1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_c_0_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5438\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => \buart.Z_rx.bitcount_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4035\,
            in2 => \_gnd_net_\,
            in3 => \N__3772\,
            lcout => \buart.Z_rx.bitcount_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_0\,
            carryout => \buart.Z_rx.bitcount_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3853\,
            in2 => \_gnd_net_\,
            in3 => \N__3769\,
            lcout => \buart.Z_rx.bitcount_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_1\,
            carryout => \buart.Z_rx.bitcount_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4122\,
            in2 => \_gnd_net_\,
            in3 => \N__3766\,
            lcout => \buart.Z_rx.bitcount_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_2\,
            carryout => \buart.Z_rx.bitcount_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNO_0_4_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101101001110"
        )
    port map (
            in0 => \N__3985\,
            in1 => \N__4177\,
            in2 => \N__3928\,
            in3 => \N__3763\,
            lcout => \buart.Z_rx.bitcount_lm_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNO_0_1_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101100110"
        )
    port map (
            in0 => \N__3754\,
            in1 => \N__4036\,
            in2 => \N__3927\,
            in3 => \N__3986\,
            lcout => \buart.Z_rx.bitcount_lm_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNO_0_3_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101100110"
        )
    port map (
            in0 => \N__4123\,
            in1 => \N__3748\,
            in2 => \N__3941\,
            in3 => \N__3988\,
            lcout => OPEN,
            ltout => \buart.Z_rx.bitcount_lm_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_3_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__4121\,
            in1 => \N__3969\,
            in2 => \N__3742\,
            in3 => \N__3923\,
            lcout => \buart__rx_bitcount_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6171\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNIMK771_4_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3850\,
            in1 => \N__4030\,
            in2 => \N__4180\,
            in3 => \N__4120\,
            lcout => OPEN,
            ltout => \buart.Z_rx.bitcount_RNIMK771Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNI9F1H1_0_0_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4078\,
            in3 => \N__5437\,
            lcout => \buart.Z_rx.idle\,
            ltout => \buart.Z_rx.idle_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.hh_RNI065O1_0_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4218\,
            in2 => \N__4066\,
            in3 => \N__4063\,
            lcout => \buart.Z_rx.startbit\,
            ltout => \buart.Z_rx.startbit_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_1_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101100001000"
        )
    port map (
            in0 => \N__4031\,
            in1 => \N__3967\,
            in2 => \N__4045\,
            in3 => \N__4042\,
            lcout => \buart__rx_bitcount_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6171\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNO_0_2_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101100110"
        )
    port map (
            in0 => \N__3851\,
            in1 => \N__3994\,
            in2 => \N__3940\,
            in3 => \N__3987\,
            lcout => OPEN,
            ltout => \buart.Z_rx.bitcount_lm_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_2_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__3854\,
            in1 => \N__3968\,
            in2 => \N__3949\,
            in3 => \N__3922\,
            lcout => \buart__rx_bitcount_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6171\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.de0.g0_13_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__6659\,
            in1 => \N__6446\,
            in2 => \N__6535\,
            in3 => \N__6576\,
            lcout => \Glue_Lab2.g0_8_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_3_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5495\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6175\,
            ce => \N__6073\,
            sr => \_gnd_net_\
        );

    \Glue_Lab2.de0.un2_de_hexplus_2_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__5101\,
            in1 => \_gnd_net_\,
            in2 => \N__6673\,
            in3 => \N__6572\,
            lcout => \Glue_Lab2.de0.un2_de_hexplusZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_6_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6660\,
            lcout => bu_rx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6175\,
            ce => \N__6073\,
            sr => \_gnd_net_\
        );

    \Glue_Lab2.de0.un1_charData_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__5100\,
            in1 => \N__4230\,
            in2 => \N__6672\,
            in3 => \N__5493\,
            lcout => \Glue_Lab2.de0.un1_charDataZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_fast_5_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5103\,
            lcout => \buart__rx_shifter_fast_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6175\,
            ce => \N__6073\,
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_7_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4219\,
            lcout => bu_rx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6175\,
            ce => \N__6073\,
            sr => \_gnd_net_\
        );

    \Glue_Lab2.gl_fsm.enOp_0_a2_4_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__5494\,
            in1 => \N__6530\,
            in2 => \N__6595\,
            in3 => \N__5102\,
            lcout => \Glue_Lab2.gl_fsm.enOp_0_a2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.de0.g0_1_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__6662\,
            in1 => \N__6578\,
            in2 => \N__6534\,
            in3 => \N__6460\,
            lcout => \Glue_Lab2.g0_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_1_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5226\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6180\,
            ce => \N__6058\,
            sr => \_gnd_net_\
        );

    \Glue_Lab2.de0.de_esc_3_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6661\,
            in1 => \N__6577\,
            in2 => \_gnd_net_\,
            in3 => \N__6461\,
            lcout => \Glue_Lab2.de0.de_escZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_0_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6462\,
            lcout => bu_rx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6180\,
            ce => \N__6058\,
            sr => \_gnd_net_\
        );

    \Glue_Lab2.gl_fsm.state_RNIQ3DV3_0_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4666\,
            in1 => \N__4330\,
            in2 => \N__4324\,
            in3 => \N__4315\,
            lcout => \Glue_Lab2.enOp\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_rst_RNI7BQG_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6450\,
            in2 => \_gnd_net_\,
            in3 => \N__6309\,
            lcout => OPEN,
            ltout => \Glue_Lab2.Gl_r1_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_Op_1_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__5977\,
            in1 => \N__6337\,
            in2 => \N__4294\,
            in3 => \N__4274\,
            lcout => \Glue_Lab2_Gl_Op_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6186\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_rst_RNI8CQG_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6310\,
            in2 => \_gnd_net_\,
            in3 => \N__5231\,
            lcout => OPEN,
            ltout => \Glue_Lab2.Gl_r1_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_Op_2_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__6311\,
            in1 => \N__4275\,
            in2 => \N__4291\,
            in3 => \N__5916\,
            lcout => \Glue_Lab2_Gl_Op_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6186\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_Op_5_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__4273\,
            in1 => \N__6313\,
            in2 => \_gnd_net_\,
            in3 => \N__5951\,
            lcout => \Glue_Lab2_Gl_Op_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6186\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.g0_1_2_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6029\,
            in1 => \N__6005\,
            in2 => \N__5982\,
            in3 => \N__5915\,
            lcout => \Lab_UT.g0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_Op_3_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111010"
        )
    port map (
            in0 => \N__6006\,
            in1 => \_gnd_net_\,
            in2 => \N__4276\,
            in3 => \N__6312\,
            lcout => \Glue_Lab2_Gl_Op_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6186\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_Op_0_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__6030\,
            in1 => \N__6336\,
            in2 => \_gnd_net_\,
            in3 => \N__4269\,
            lcout => \Glue_Lab2_Gl_Op_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6186\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_tx_data_2_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__4614\,
            in1 => \N__5032\,
            in2 => \_gnd_net_\,
            in3 => \N__5236\,
            lcout => \Gl_tx_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6190\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.gl_fsm.state_RNIIM7B_1_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4689\,
            in2 => \_gnd_net_\,
            in3 => \N__6674\,
            lcout => \Glue_Lab2.gl_fsm.enOp_0_a2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_Op_RNIDA8P_2_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6001\,
            in2 => \_gnd_net_\,
            in3 => \N__5914\,
            lcout => OPEN,
            ltout => \Glue_Lab2.Gl_subtract_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_Op_RNIFO4V1_0_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5952\,
            in1 => \N__5981\,
            in2 => \N__4657\,
            in3 => \N__6025\,
            lcout => \Gl_subtract\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.S_0_s_ac0_5_d_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000010000000"
        )
    port map (
            in0 => \N__5862\,
            in1 => \N__4654\,
            in2 => \N__4645\,
            in3 => \N__5780\,
            lcout => \Lab_UT.S_0_s_ac0_5_dZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.S_m_am_2_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__5779\,
            in1 => \N__5861\,
            in2 => \_gnd_net_\,
            in3 => \N__4641\,
            lcout => OPEN,
            ltout => \Lab_UT.S_m_amZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.S_m_ns_2_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4717\,
            in2 => \N__4624\,
            in3 => \N__5557\,
            lcout => led_c_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.S_m_bm_1_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001110011100"
        )
    port map (
            in0 => \N__4597\,
            in1 => \N__4548\,
            in2 => \N__4488\,
            in3 => \N__4420\,
            lcout => OPEN,
            ltout => \Lab_UT.S_m_bmZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.S_m_ns_1_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4351\,
            in2 => \N__4345\,
            in3 => \N__5558\,
            lcout => led_c_1,
            ltout => \led_c_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_tx_data_1_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6470\,
            in2 => \N__4765\,
            in3 => \N__5033\,
            lcout => \Gl_tx_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6193\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.S_m_bm_2_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__4750\,
            in1 => \N__4735\,
            in2 => \_gnd_net_\,
            in3 => \N__4723\,
            lcout => \Lab_UT.S_m_bmZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNI1O14_1_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4839\,
            in2 => \_gnd_net_\,
            in3 => \N__4817\,
            lcout => \buart.Z_tx.Z_baudgen.un2_counter_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_0_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4818\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6182\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_1_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__4819\,
            in1 => \_gnd_net_\,
            in2 => \N__4843\,
            in3 => \_gnd_net_\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6182\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_4_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__4888\,
            in1 => \N__6820\,
            in2 => \N__6886\,
            in3 => \N__6908\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6177\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNIQJ4A_4_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6907\,
            in1 => \N__4887\,
            in2 => \N__6823\,
            in3 => \N__6881\,
            lcout => \buart.Z_tx.Z_baudgen.un2_counter_c5\,
            ltout => \buart.Z_tx.Z_baudgen.un2_counter_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_5_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001011010"
        )
    port map (
            in0 => \N__4871\,
            in1 => \_gnd_net_\,
            in2 => \N__4711\,
            in3 => \N__6855\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6177\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNINP26_6_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__4853\,
            in1 => \N__4837\,
            in2 => \_gnd_net_\,
            in3 => \N__4815\,
            lcout => \buart.Z_tx.Z_baudgen.un1_bitcount_c2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_6_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__4872\,
            in1 => \N__4855\,
            in2 => \N__4708\,
            in3 => \N__6856\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6177\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNIES38_0_4_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__6906\,
            in1 => \N__4886\,
            in2 => \N__6822\,
            in3 => \N__4870\,
            lcout => \buart.Z_tx.Z_baudgen.counter_RNIES38_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNIES38_4_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__4885\,
            in1 => \N__6813\,
            in2 => \N__4873\,
            in3 => \N__6905\,
            lcout => OPEN,
            ltout => \buart.Z_tx.Z_baudgen.ser_clk_sx_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNI5M6E_6_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__4854\,
            in1 => \N__4838\,
            in2 => \N__4822\,
            in3 => \N__4816\,
            lcout => \buart.Z_tx.ser_clk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNIBADL_1_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4959\,
            in2 => \_gnd_net_\,
            in3 => \N__4919\,
            lcout => OPEN,
            ltout => \buart.Z_tx.bitcount_RNIBADLZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNIVE1P1_4_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000100010"
        )
    port map (
            in0 => \N__4798\,
            in1 => \N__4792\,
            in2 => \N__4786\,
            in3 => \N__4774\,
            lcout => \buart.Z_tx.counter_RNIVE1P1_4\,
            ltout => \buart.Z_tx.counter_RNIVE1P1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_2_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__6786\,
            in1 => \N__5068\,
            in2 => \N__4783\,
            in3 => \N__4780\,
            lcout => \buart.Z_tx.bitcountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6172\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNO_0_2_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__4921\,
            in1 => \N__4961\,
            in2 => \_gnd_net_\,
            in3 => \N__6848\,
            lcout => \buart.Z_tx.un1_bitcount_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNIFEDL_3_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5052\,
            in2 => \_gnd_net_\,
            in3 => \N__5066\,
            lcout => \buart.Z_tx.uart_busy_0_0\,
            ltout => \buart.Z_tx.uart_busy_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNIQL5G1_1_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__4920\,
            in1 => \N__6785\,
            in2 => \N__4768\,
            in3 => \N__4960\,
            lcout => \buart.Z_tx.un1_uart_wr_i_0_i_sx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNO_0_3_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__6849\,
            in1 => \N__4922\,
            in2 => \N__4966\,
            in3 => \N__5067\,
            lcout => OPEN,
            ltout => \buart.Z_tx.un1_bitcount_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_3_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110111011110"
        )
    port map (
            in0 => \N__5053\,
            in1 => \N__6787\,
            in2 => \N__5056\,
            in3 => \N__4939\,
            lcout => \buart.Z_tx.bitcountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6172\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNIV8N32_1_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__6859\,
            in1 => \N__6761\,
            in2 => \_gnd_net_\,
            in3 => \N__5044\,
            lcout => \buart.Z_tx.un1_uart_wr_i_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_tx_data_rdy_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__6202\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5038\,
            lcout => \Gl_tx_data_rdy\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6176\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNO_0_1_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4923\,
            in2 => \_gnd_net_\,
            in3 => \N__6858\,
            lcout => OPEN,
            ltout => \buart.Z_tx.un1_bitcount_c1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_1_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110111011110"
        )
    port map (
            in0 => \N__4938\,
            in1 => \N__6763\,
            in2 => \N__4969\,
            in3 => \N__4965\,
            lcout => \buart.Z_tx.bitcountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6176\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_0_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6762\,
            in1 => \N__4924\,
            in2 => \_gnd_net_\,
            in3 => \N__4937\,
            lcout => \buart.Z_tx.bitcountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6176\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.de0.de_esc_4_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__5487\,
            in1 => \N__6505\,
            in2 => \N__5129\,
            in3 => \N__5175\,
            lcout => \Glue_Lab2.de0.de_escZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.de0.g0_10_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5118\,
            in2 => \_gnd_net_\,
            in3 => \N__5489\,
            lcout => OPEN,
            ltout => \Glue_Lab2.de0.g0_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.de0.g0_3_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__5454\,
            in1 => \N__5177\,
            in2 => \N__5527\,
            in3 => \N__5385\,
            lcout => OPEN,
            ltout => \Glue_Lab2.g0_9_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.reset_count_RNO_0_1_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__5303\,
            in1 => \N__6388\,
            in2 => \N__5524\,
            in3 => \N__5521\,
            lcout => \Glue_Lab2.reset_counte_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_4_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6506\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6181\,
            ce => \N__6072\,
            sr => \_gnd_net_\
        );

    \Glue_Lab2.de0.g0_5_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5119\,
            in2 => \_gnd_net_\,
            in3 => \N__5488\,
            lcout => OPEN,
            ltout => \Glue_Lab2.de0.g0Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.de0.g0_9_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__5455\,
            in1 => \N__5176\,
            in2 => \N__5392\,
            in3 => \N__5384\,
            lcout => OPEN,
            ltout => \Glue_Lab2.g0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.reset_count_RNO_0_3_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__5304\,
            in1 => \N__6685\,
            in2 => \N__5260\,
            in3 => \N__5257\,
            lcout => \Glue_Lab2.reset_counte_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_2_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6613\,
            lcout => bu_rx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6187\,
            ce => \N__6071\,
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_5_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5131\,
            lcout => bu_rx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6187\,
            ce => \N__6071\,
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_fast_4_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6519\,
            lcout => \buart__rx_shifter_fast_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6187\,
            ce => \N__6071\,
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_tx_data_RNO_1_5_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6031\,
            in2 => \_gnd_net_\,
            in3 => \N__6007\,
            lcout => OPEN,
            ltout => \Glue_Lab2.g0_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.Gl_tx_data_RNO_0_5_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__5983\,
            in1 => \N__5953\,
            in2 => \N__5923\,
            in3 => \N__5920\,
            lcout => \Glue_Lab2.Gl_subtract_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.S_0_s_ac0_5_0_0_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010000000"
        )
    port map (
            in0 => \N__5883\,
            in1 => \N__5814\,
            in2 => \N__5662\,
            in3 => \N__5733\,
            lcout => \Lab_UT.S_0_s_ac0_5_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.S_1_c3_c_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__5884\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5815\,
            lcout => OPEN,
            ltout => \Lab_UT.S_1_c3_cZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.S_1_c4_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011101010"
        )
    port map (
            in0 => \N__5734\,
            in1 => \N__5677\,
            in2 => \N__5665\,
            in3 => \N__5660\,
            lcout => OPEN,
            ltout => \Lab_UT.C_out41_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.L2_led_1_4_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111101110"
        )
    port map (
            in0 => \N__5593\,
            in1 => \N__5587\,
            in2 => \N__5575\,
            in3 => \N__5572\,
            lcout => led_c_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_2_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6877\,
            in2 => \_gnd_net_\,
            in3 => \N__6909\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6184\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_3_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__6910\,
            in1 => \N__6821\,
            in2 => \N__6885\,
            in3 => \N__6857\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6184\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_8_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6764\,
            lcout => \buart.Z_tx.shifterZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6183\,
            ce => \N__6701\,
            sr => \_gnd_net_\
        );

    \Glue_Lab2.de0.g0_8_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__6675\,
            in1 => \N__6596\,
            in2 => \N__6529\,
            in3 => \N__6472\,
            lcout => \Glue_Lab2.g0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.sDelay.delayReg_3_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__6307\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6373\,
            lcout => \Lab_UT.sDelay.delayRegZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6191\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Glue_Lab2.de0.g0_6_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__6679\,
            in1 => \N__6612\,
            in2 => \N__6528\,
            in3 => \N__6473\,
            lcout => \Glue_Lab2.g0_8_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.sDelay.delayReg_2_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__6306\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6382\,
            lcout => \Lab_UT.sDelay.delayRegZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6191\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.sDelay.delayReg_4_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6367\,
            in2 => \_gnd_net_\,
            in3 => \N__6308\,
            lcout => \L2_adder_rdy\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6191\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
