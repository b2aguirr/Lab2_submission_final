// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     May 1 2019 17:42:51

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "latticehx1k" view "INTERFACE"

module latticehx1k (
    led,
    to_ir,
    test2,
    sd,
    test1,
    o_serial_data,
    from_pc,
    test3,
    clk_in);

    output [4:0] led;
    output to_ir;
    output test2;
    output sd;
    output test1;
    output o_serial_data;
    input from_pc;
    output test3;
    input clk_in;

    wire N__7037;
    wire N__7036;
    wire N__7035;
    wire N__7028;
    wire N__7027;
    wire N__7026;
    wire N__7019;
    wire N__7018;
    wire N__7017;
    wire N__7010;
    wire N__7009;
    wire N__7008;
    wire N__7001;
    wire N__7000;
    wire N__6999;
    wire N__6992;
    wire N__6991;
    wire N__6990;
    wire N__6983;
    wire N__6982;
    wire N__6981;
    wire N__6974;
    wire N__6973;
    wire N__6972;
    wire N__6965;
    wire N__6964;
    wire N__6963;
    wire N__6956;
    wire N__6955;
    wire N__6954;
    wire N__6947;
    wire N__6946;
    wire N__6945;
    wire N__6938;
    wire N__6937;
    wire N__6936;
    wire N__6929;
    wire N__6928;
    wire N__6927;
    wire N__6910;
    wire N__6909;
    wire N__6908;
    wire N__6907;
    wire N__6906;
    wire N__6905;
    wire N__6900;
    wire N__6891;
    wire N__6886;
    wire N__6885;
    wire N__6882;
    wire N__6881;
    wire N__6878;
    wire N__6877;
    wire N__6872;
    wire N__6867;
    wire N__6864;
    wire N__6859;
    wire N__6858;
    wire N__6857;
    wire N__6856;
    wire N__6855;
    wire N__6850;
    wire N__6849;
    wire N__6848;
    wire N__6845;
    wire N__6840;
    wire N__6837;
    wire N__6832;
    wire N__6823;
    wire N__6822;
    wire N__6821;
    wire N__6820;
    wire N__6817;
    wire N__6814;
    wire N__6813;
    wire N__6810;
    wire N__6801;
    wire N__6796;
    wire N__6795;
    wire N__6794;
    wire N__6793;
    wire N__6792;
    wire N__6791;
    wire N__6790;
    wire N__6789;
    wire N__6788;
    wire N__6787;
    wire N__6786;
    wire N__6785;
    wire N__6782;
    wire N__6765;
    wire N__6764;
    wire N__6763;
    wire N__6762;
    wire N__6761;
    wire N__6754;
    wire N__6749;
    wire N__6746;
    wire N__6739;
    wire N__6736;
    wire N__6727;
    wire N__6724;
    wire N__6721;
    wire N__6718;
    wire N__6715;
    wire N__6712;
    wire N__6711;
    wire N__6708;
    wire N__6705;
    wire N__6702;
    wire N__6701;
    wire N__6698;
    wire N__6695;
    wire N__6692;
    wire N__6685;
    wire N__6682;
    wire N__6679;
    wire N__6676;
    wire N__6675;
    wire N__6674;
    wire N__6673;
    wire N__6672;
    wire N__6669;
    wire N__6666;
    wire N__6663;
    wire N__6662;
    wire N__6661;
    wire N__6660;
    wire N__6659;
    wire N__6656;
    wire N__6653;
    wire N__6650;
    wire N__6647;
    wire N__6644;
    wire N__6639;
    wire N__6630;
    wire N__6619;
    wire N__6616;
    wire N__6615;
    wire N__6614;
    wire N__6613;
    wire N__6612;
    wire N__6609;
    wire N__6606;
    wire N__6603;
    wire N__6600;
    wire N__6597;
    wire N__6596;
    wire N__6595;
    wire N__6590;
    wire N__6587;
    wire N__6582;
    wire N__6579;
    wire N__6578;
    wire N__6577;
    wire N__6576;
    wire N__6573;
    wire N__6572;
    wire N__6569;
    wire N__6566;
    wire N__6563;
    wire N__6560;
    wire N__6555;
    wire N__6548;
    wire N__6535;
    wire N__6534;
    wire N__6531;
    wire N__6530;
    wire N__6529;
    wire N__6528;
    wire N__6525;
    wire N__6520;
    wire N__6519;
    wire N__6516;
    wire N__6513;
    wire N__6510;
    wire N__6507;
    wire N__6506;
    wire N__6505;
    wire N__6502;
    wire N__6499;
    wire N__6496;
    wire N__6491;
    wire N__6486;
    wire N__6475;
    wire N__6474;
    wire N__6473;
    wire N__6472;
    wire N__6471;
    wire N__6470;
    wire N__6469;
    wire N__6466;
    wire N__6463;
    wire N__6462;
    wire N__6461;
    wire N__6460;
    wire N__6457;
    wire N__6454;
    wire N__6451;
    wire N__6450;
    wire N__6447;
    wire N__6446;
    wire N__6443;
    wire N__6438;
    wire N__6431;
    wire N__6428;
    wire N__6425;
    wire N__6422;
    wire N__6419;
    wire N__6416;
    wire N__6413;
    wire N__6410;
    wire N__6399;
    wire N__6388;
    wire N__6385;
    wire N__6382;
    wire N__6379;
    wire N__6376;
    wire N__6373;
    wire N__6370;
    wire N__6367;
    wire N__6364;
    wire N__6361;
    wire N__6360;
    wire N__6359;
    wire N__6358;
    wire N__6357;
    wire N__6356;
    wire N__6355;
    wire N__6354;
    wire N__6353;
    wire N__6352;
    wire N__6349;
    wire N__6348;
    wire N__6345;
    wire N__6344;
    wire N__6343;
    wire N__6340;
    wire N__6339;
    wire N__6338;
    wire N__6337;
    wire N__6336;
    wire N__6333;
    wire N__6324;
    wire N__6319;
    wire N__6314;
    wire N__6313;
    wire N__6312;
    wire N__6311;
    wire N__6310;
    wire N__6309;
    wire N__6308;
    wire N__6307;
    wire N__6306;
    wire N__6301;
    wire N__6292;
    wire N__6291;
    wire N__6286;
    wire N__6277;
    wire N__6266;
    wire N__6259;
    wire N__6256;
    wire N__6253;
    wire N__6250;
    wire N__6249;
    wire N__6248;
    wire N__6247;
    wire N__6246;
    wire N__6239;
    wire N__6236;
    wire N__6229;
    wire N__6226;
    wire N__6223;
    wire N__6218;
    wire N__6215;
    wire N__6202;
    wire N__6199;
    wire N__6196;
    wire N__6193;
    wire N__6192;
    wire N__6191;
    wire N__6190;
    wire N__6189;
    wire N__6188;
    wire N__6187;
    wire N__6186;
    wire N__6185;
    wire N__6184;
    wire N__6183;
    wire N__6182;
    wire N__6181;
    wire N__6180;
    wire N__6179;
    wire N__6178;
    wire N__6177;
    wire N__6176;
    wire N__6175;
    wire N__6174;
    wire N__6173;
    wire N__6172;
    wire N__6171;
    wire N__6170;
    wire N__6169;
    wire N__6168;
    wire N__6167;
    wire N__6166;
    wire N__6165;
    wire N__6164;
    wire N__6163;
    wire N__6162;
    wire N__6097;
    wire N__6094;
    wire N__6091;
    wire N__6090;
    wire N__6087;
    wire N__6084;
    wire N__6081;
    wire N__6076;
    wire N__6073;
    wire N__6072;
    wire N__6071;
    wire N__6068;
    wire N__6065;
    wire N__6062;
    wire N__6059;
    wire N__6058;
    wire N__6055;
    wire N__6052;
    wire N__6049;
    wire N__6046;
    wire N__6041;
    wire N__6036;
    wire N__6031;
    wire N__6030;
    wire N__6029;
    wire N__6026;
    wire N__6025;
    wire N__6020;
    wire N__6017;
    wire N__6014;
    wire N__6007;
    wire N__6006;
    wire N__6005;
    wire N__6002;
    wire N__6001;
    wire N__5996;
    wire N__5993;
    wire N__5990;
    wire N__5983;
    wire N__5982;
    wire N__5981;
    wire N__5978;
    wire N__5977;
    wire N__5974;
    wire N__5971;
    wire N__5968;
    wire N__5963;
    wire N__5960;
    wire N__5953;
    wire N__5952;
    wire N__5951;
    wire N__5950;
    wire N__5947;
    wire N__5944;
    wire N__5941;
    wire N__5938;
    wire N__5935;
    wire N__5932;
    wire N__5923;
    wire N__5920;
    wire N__5917;
    wire N__5916;
    wire N__5915;
    wire N__5914;
    wire N__5911;
    wire N__5906;
    wire N__5903;
    wire N__5896;
    wire N__5893;
    wire N__5890;
    wire N__5887;
    wire N__5884;
    wire N__5883;
    wire N__5882;
    wire N__5877;
    wire N__5874;
    wire N__5873;
    wire N__5872;
    wire N__5871;
    wire N__5868;
    wire N__5865;
    wire N__5864;
    wire N__5863;
    wire N__5862;
    wire N__5861;
    wire N__5860;
    wire N__5857;
    wire N__5854;
    wire N__5851;
    wire N__5846;
    wire N__5841;
    wire N__5836;
    wire N__5833;
    wire N__5830;
    wire N__5815;
    wire N__5814;
    wire N__5813;
    wire N__5812;
    wire N__5811;
    wire N__5806;
    wire N__5805;
    wire N__5802;
    wire N__5801;
    wire N__5800;
    wire N__5797;
    wire N__5794;
    wire N__5791;
    wire N__5788;
    wire N__5785;
    wire N__5784;
    wire N__5781;
    wire N__5780;
    wire N__5779;
    wire N__5776;
    wire N__5773;
    wire N__5770;
    wire N__5763;
    wire N__5760;
    wire N__5757;
    wire N__5752;
    wire N__5749;
    wire N__5734;
    wire N__5733;
    wire N__5728;
    wire N__5725;
    wire N__5724;
    wire N__5723;
    wire N__5722;
    wire N__5721;
    wire N__5720;
    wire N__5719;
    wire N__5718;
    wire N__5717;
    wire N__5716;
    wire N__5715;
    wire N__5712;
    wire N__5707;
    wire N__5702;
    wire N__5695;
    wire N__5688;
    wire N__5677;
    wire N__5674;
    wire N__5671;
    wire N__5668;
    wire N__5665;
    wire N__5662;
    wire N__5661;
    wire N__5660;
    wire N__5657;
    wire N__5656;
    wire N__5653;
    wire N__5652;
    wire N__5651;
    wire N__5646;
    wire N__5643;
    wire N__5642;
    wire N__5641;
    wire N__5634;
    wire N__5633;
    wire N__5632;
    wire N__5631;
    wire N__5630;
    wire N__5627;
    wire N__5620;
    wire N__5617;
    wire N__5612;
    wire N__5607;
    wire N__5602;
    wire N__5593;
    wire N__5590;
    wire N__5587;
    wire N__5584;
    wire N__5581;
    wire N__5578;
    wire N__5575;
    wire N__5572;
    wire N__5571;
    wire N__5568;
    wire N__5565;
    wire N__5562;
    wire N__5559;
    wire N__5558;
    wire N__5557;
    wire N__5552;
    wire N__5547;
    wire N__5542;
    wire N__5539;
    wire N__5536;
    wire N__5533;
    wire N__5530;
    wire N__5527;
    wire N__5524;
    wire N__5521;
    wire N__5518;
    wire N__5515;
    wire N__5512;
    wire N__5509;
    wire N__5506;
    wire N__5503;
    wire N__5500;
    wire N__5499;
    wire N__5496;
    wire N__5495;
    wire N__5494;
    wire N__5493;
    wire N__5490;
    wire N__5489;
    wire N__5488;
    wire N__5487;
    wire N__5484;
    wire N__5477;
    wire N__5474;
    wire N__5467;
    wire N__5462;
    wire N__5455;
    wire N__5454;
    wire N__5453;
    wire N__5448;
    wire N__5447;
    wire N__5444;
    wire N__5443;
    wire N__5440;
    wire N__5439;
    wire N__5438;
    wire N__5437;
    wire N__5436;
    wire N__5435;
    wire N__5432;
    wire N__5429;
    wire N__5426;
    wire N__5423;
    wire N__5420;
    wire N__5417;
    wire N__5414;
    wire N__5409;
    wire N__5392;
    wire N__5389;
    wire N__5388;
    wire N__5387;
    wire N__5386;
    wire N__5385;
    wire N__5384;
    wire N__5383;
    wire N__5382;
    wire N__5377;
    wire N__5374;
    wire N__5371;
    wire N__5366;
    wire N__5363;
    wire N__5360;
    wire N__5357;
    wire N__5356;
    wire N__5355;
    wire N__5352;
    wire N__5349;
    wire N__5346;
    wire N__5345;
    wire N__5344;
    wire N__5341;
    wire N__5336;
    wire N__5331;
    wire N__5328;
    wire N__5323;
    wire N__5318;
    wire N__5305;
    wire N__5304;
    wire N__5303;
    wire N__5300;
    wire N__5295;
    wire N__5294;
    wire N__5293;
    wire N__5292;
    wire N__5289;
    wire N__5286;
    wire N__5283;
    wire N__5280;
    wire N__5277;
    wire N__5274;
    wire N__5269;
    wire N__5260;
    wire N__5257;
    wire N__5254;
    wire N__5251;
    wire N__5248;
    wire N__5245;
    wire N__5242;
    wire N__5239;
    wire N__5236;
    wire N__5235;
    wire N__5234;
    wire N__5233;
    wire N__5232;
    wire N__5231;
    wire N__5230;
    wire N__5229;
    wire N__5228;
    wire N__5227;
    wire N__5226;
    wire N__5223;
    wire N__5220;
    wire N__5213;
    wire N__5210;
    wire N__5207;
    wire N__5204;
    wire N__5201;
    wire N__5198;
    wire N__5197;
    wire N__5196;
    wire N__5193;
    wire N__5184;
    wire N__5181;
    wire N__5178;
    wire N__5177;
    wire N__5176;
    wire N__5175;
    wire N__5170;
    wire N__5167;
    wire N__5164;
    wire N__5157;
    wire N__5154;
    wire N__5147;
    wire N__5140;
    wire N__5131;
    wire N__5130;
    wire N__5129;
    wire N__5126;
    wire N__5123;
    wire N__5120;
    wire N__5119;
    wire N__5118;
    wire N__5115;
    wire N__5112;
    wire N__5105;
    wire N__5104;
    wire N__5103;
    wire N__5102;
    wire N__5101;
    wire N__5100;
    wire N__5099;
    wire N__5092;
    wire N__5089;
    wire N__5080;
    wire N__5077;
    wire N__5068;
    wire N__5067;
    wire N__5066;
    wire N__5059;
    wire N__5056;
    wire N__5053;
    wire N__5052;
    wire N__5047;
    wire N__5044;
    wire N__5041;
    wire N__5038;
    wire N__5037;
    wire N__5034;
    wire N__5033;
    wire N__5032;
    wire N__5031;
    wire N__5028;
    wire N__5025;
    wire N__5022;
    wire N__5019;
    wire N__5018;
    wire N__5017;
    wire N__5016;
    wire N__5011;
    wire N__5010;
    wire N__5009;
    wire N__5008;
    wire N__5005;
    wire N__5000;
    wire N__4995;
    wire N__4992;
    wire N__4989;
    wire N__4982;
    wire N__4969;
    wire N__4966;
    wire N__4965;
    wire N__4962;
    wire N__4961;
    wire N__4960;
    wire N__4959;
    wire N__4956;
    wire N__4949;
    wire N__4946;
    wire N__4939;
    wire N__4938;
    wire N__4937;
    wire N__4934;
    wire N__4929;
    wire N__4924;
    wire N__4923;
    wire N__4922;
    wire N__4921;
    wire N__4920;
    wire N__4919;
    wire N__4914;
    wire N__4905;
    wire N__4900;
    wire N__4897;
    wire N__4894;
    wire N__4891;
    wire N__4888;
    wire N__4887;
    wire N__4886;
    wire N__4885;
    wire N__4876;
    wire N__4873;
    wire N__4872;
    wire N__4871;
    wire N__4870;
    wire N__4867;
    wire N__4858;
    wire N__4855;
    wire N__4854;
    wire N__4853;
    wire N__4846;
    wire N__4843;
    wire N__4840;
    wire N__4839;
    wire N__4838;
    wire N__4837;
    wire N__4832;
    wire N__4827;
    wire N__4822;
    wire N__4819;
    wire N__4818;
    wire N__4817;
    wire N__4816;
    wire N__4815;
    wire N__4808;
    wire N__4803;
    wire N__4798;
    wire N__4795;
    wire N__4792;
    wire N__4789;
    wire N__4786;
    wire N__4783;
    wire N__4780;
    wire N__4777;
    wire N__4774;
    wire N__4771;
    wire N__4768;
    wire N__4765;
    wire N__4762;
    wire N__4759;
    wire N__4756;
    wire N__4753;
    wire N__4750;
    wire N__4747;
    wire N__4746;
    wire N__4743;
    wire N__4740;
    wire N__4735;
    wire N__4734;
    wire N__4731;
    wire N__4728;
    wire N__4723;
    wire N__4720;
    wire N__4717;
    wire N__4714;
    wire N__4711;
    wire N__4708;
    wire N__4705;
    wire N__4702;
    wire N__4699;
    wire N__4698;
    wire N__4697;
    wire N__4696;
    wire N__4695;
    wire N__4690;
    wire N__4689;
    wire N__4686;
    wire N__4681;
    wire N__4678;
    wire N__4675;
    wire N__4666;
    wire N__4663;
    wire N__4660;
    wire N__4657;
    wire N__4654;
    wire N__4651;
    wire N__4648;
    wire N__4645;
    wire N__4642;
    wire N__4641;
    wire N__4636;
    wire N__4635;
    wire N__4632;
    wire N__4629;
    wire N__4624;
    wire N__4621;
    wire N__4618;
    wire N__4615;
    wire N__4614;
    wire N__4611;
    wire N__4608;
    wire N__4603;
    wire N__4602;
    wire N__4601;
    wire N__4598;
    wire N__4597;
    wire N__4596;
    wire N__4595;
    wire N__4594;
    wire N__4591;
    wire N__4590;
    wire N__4587;
    wire N__4584;
    wire N__4581;
    wire N__4578;
    wire N__4569;
    wire N__4558;
    wire N__4557;
    wire N__4556;
    wire N__4553;
    wire N__4552;
    wire N__4551;
    wire N__4550;
    wire N__4549;
    wire N__4548;
    wire N__4547;
    wire N__4546;
    wire N__4543;
    wire N__4532;
    wire N__4529;
    wire N__4528;
    wire N__4527;
    wire N__4526;
    wire N__4523;
    wire N__4520;
    wire N__4515;
    wire N__4510;
    wire N__4505;
    wire N__4502;
    wire N__4489;
    wire N__4488;
    wire N__4487;
    wire N__4486;
    wire N__4485;
    wire N__4482;
    wire N__4479;
    wire N__4478;
    wire N__4475;
    wire N__4474;
    wire N__4471;
    wire N__4468;
    wire N__4465;
    wire N__4462;
    wire N__4453;
    wire N__4450;
    wire N__4449;
    wire N__4444;
    wire N__4441;
    wire N__4438;
    wire N__4435;
    wire N__4432;
    wire N__4429;
    wire N__4420;
    wire N__4417;
    wire N__4416;
    wire N__4415;
    wire N__4414;
    wire N__4411;
    wire N__4406;
    wire N__4403;
    wire N__4402;
    wire N__4401;
    wire N__4400;
    wire N__4399;
    wire N__4398;
    wire N__4397;
    wire N__4396;
    wire N__4395;
    wire N__4394;
    wire N__4391;
    wire N__4388;
    wire N__4385;
    wire N__4374;
    wire N__4367;
    wire N__4364;
    wire N__4351;
    wire N__4348;
    wire N__4345;
    wire N__4342;
    wire N__4339;
    wire N__4336;
    wire N__4333;
    wire N__4330;
    wire N__4327;
    wire N__4324;
    wire N__4321;
    wire N__4318;
    wire N__4315;
    wire N__4314;
    wire N__4313;
    wire N__4312;
    wire N__4309;
    wire N__4304;
    wire N__4301;
    wire N__4294;
    wire N__4291;
    wire N__4288;
    wire N__4285;
    wire N__4282;
    wire N__4279;
    wire N__4276;
    wire N__4275;
    wire N__4274;
    wire N__4273;
    wire N__4270;
    wire N__4269;
    wire N__4268;
    wire N__4257;
    wire N__4254;
    wire N__4249;
    wire N__4246;
    wire N__4243;
    wire N__4240;
    wire N__4237;
    wire N__4234;
    wire N__4231;
    wire N__4230;
    wire N__4227;
    wire N__4224;
    wire N__4219;
    wire N__4218;
    wire N__4215;
    wire N__4212;
    wire N__4209;
    wire N__4206;
    wire N__4201;
    wire N__4198;
    wire N__4195;
    wire N__4192;
    wire N__4189;
    wire N__4186;
    wire N__4183;
    wire N__4182;
    wire N__4181;
    wire N__4180;
    wire N__4179;
    wire N__4178;
    wire N__4177;
    wire N__4174;
    wire N__4171;
    wire N__4168;
    wire N__4165;
    wire N__4164;
    wire N__4161;
    wire N__4160;
    wire N__4157;
    wire N__4154;
    wire N__4151;
    wire N__4146;
    wire N__4143;
    wire N__4136;
    wire N__4123;
    wire N__4122;
    wire N__4121;
    wire N__4120;
    wire N__4119;
    wire N__4118;
    wire N__4117;
    wire N__4116;
    wire N__4115;
    wire N__4114;
    wire N__4111;
    wire N__4108;
    wire N__4103;
    wire N__4096;
    wire N__4089;
    wire N__4078;
    wire N__4075;
    wire N__4074;
    wire N__4069;
    wire N__4066;
    wire N__4063;
    wire N__4060;
    wire N__4059;
    wire N__4056;
    wire N__4053;
    wire N__4050;
    wire N__4045;
    wire N__4042;
    wire N__4039;
    wire N__4036;
    wire N__4035;
    wire N__4034;
    wire N__4033;
    wire N__4032;
    wire N__4031;
    wire N__4030;
    wire N__4029;
    wire N__4028;
    wire N__4027;
    wire N__4022;
    wire N__4015;
    wire N__4010;
    wire N__4003;
    wire N__3994;
    wire N__3991;
    wire N__3988;
    wire N__3987;
    wire N__3986;
    wire N__3985;
    wire N__3980;
    wire N__3975;
    wire N__3970;
    wire N__3969;
    wire N__3968;
    wire N__3967;
    wire N__3964;
    wire N__3957;
    wire N__3954;
    wire N__3949;
    wire N__3946;
    wire N__3945;
    wire N__3944;
    wire N__3943;
    wire N__3942;
    wire N__3941;
    wire N__3940;
    wire N__3937;
    wire N__3934;
    wire N__3929;
    wire N__3928;
    wire N__3927;
    wire N__3924;
    wire N__3923;
    wire N__3922;
    wire N__3919;
    wire N__3916;
    wire N__3909;
    wire N__3908;
    wire N__3907;
    wire N__3906;
    wire N__3905;
    wire N__3902;
    wire N__3899;
    wire N__3896;
    wire N__3887;
    wire N__3884;
    wire N__3875;
    wire N__3872;
    wire N__3869;
    wire N__3856;
    wire N__3855;
    wire N__3854;
    wire N__3853;
    wire N__3852;
    wire N__3851;
    wire N__3850;
    wire N__3849;
    wire N__3848;
    wire N__3845;
    wire N__3844;
    wire N__3841;
    wire N__3838;
    wire N__3835;
    wire N__3832;
    wire N__3827;
    wire N__3822;
    wire N__3815;
    wire N__3802;
    wire N__3799;
    wire N__3796;
    wire N__3793;
    wire N__3790;
    wire N__3787;
    wire N__3784;
    wire N__3781;
    wire N__3778;
    wire N__3775;
    wire N__3772;
    wire N__3769;
    wire N__3766;
    wire N__3763;
    wire N__3760;
    wire N__3757;
    wire N__3754;
    wire N__3751;
    wire N__3748;
    wire N__3745;
    wire N__3742;
    wire N__3739;
    wire N__3736;
    wire N__3733;
    wire N__3730;
    wire N__3727;
    wire N__3726;
    wire N__3725;
    wire N__3724;
    wire N__3721;
    wire N__3718;
    wire N__3713;
    wire N__3706;
    wire N__3705;
    wire N__3704;
    wire N__3703;
    wire N__3700;
    wire N__3697;
    wire N__3690;
    wire N__3687;
    wire N__3684;
    wire N__3679;
    wire N__3676;
    wire N__3673;
    wire N__3672;
    wire N__3669;
    wire N__3668;
    wire N__3665;
    wire N__3662;
    wire N__3659;
    wire N__3656;
    wire N__3653;
    wire N__3650;
    wire N__3647;
    wire N__3642;
    wire N__3637;
    wire N__3634;
    wire N__3631;
    wire N__3628;
    wire N__3627;
    wire N__3624;
    wire N__3621;
    wire N__3616;
    wire N__3613;
    wire N__3610;
    wire N__3607;
    wire N__3604;
    wire N__3601;
    wire N__3598;
    wire N__3595;
    wire N__3592;
    wire N__3589;
    wire N__3586;
    wire N__3583;
    wire N__3580;
    wire N__3579;
    wire N__3576;
    wire N__3573;
    wire N__3572;
    wire N__3567;
    wire N__3564;
    wire N__3559;
    wire N__3558;
    wire N__3557;
    wire N__3552;
    wire N__3549;
    wire N__3546;
    wire N__3543;
    wire N__3538;
    wire N__3535;
    wire N__3534;
    wire N__3533;
    wire N__3528;
    wire N__3527;
    wire N__3526;
    wire N__3523;
    wire N__3522;
    wire N__3519;
    wire N__3516;
    wire N__3513;
    wire N__3508;
    wire N__3503;
    wire N__3496;
    wire N__3493;
    wire N__3490;
    wire N__3487;
    wire N__3484;
    wire N__3481;
    wire N__3478;
    wire N__3475;
    wire N__3472;
    wire N__3469;
    wire N__3466;
    wire N__3463;
    wire N__3462;
    wire N__3459;
    wire N__3456;
    wire N__3451;
    wire N__3448;
    wire N__3447;
    wire N__3446;
    wire N__3445;
    wire N__3444;
    wire N__3443;
    wire N__3440;
    wire N__3437;
    wire N__3434;
    wire N__3427;
    wire N__3424;
    wire N__3421;
    wire N__3412;
    wire N__3409;
    wire N__3408;
    wire N__3407;
    wire N__3404;
    wire N__3401;
    wire N__3398;
    wire N__3391;
    wire N__3390;
    wire N__3387;
    wire N__3384;
    wire N__3381;
    wire N__3376;
    wire N__3375;
    wire N__3374;
    wire N__3373;
    wire N__3370;
    wire N__3367;
    wire N__3362;
    wire N__3359;
    wire N__3352;
    wire N__3349;
    wire N__3346;
    wire N__3343;
    wire N__3340;
    wire N__3337;
    wire N__3334;
    wire N__3331;
    wire N__3328;
    wire N__3325;
    wire N__3322;
    wire N__3321;
    wire N__3320;
    wire N__3319;
    wire N__3318;
    wire N__3317;
    wire N__3312;
    wire N__3307;
    wire N__3304;
    wire N__3301;
    wire N__3292;
    wire N__3291;
    wire N__3288;
    wire N__3285;
    wire N__3284;
    wire N__3283;
    wire N__3280;
    wire N__3277;
    wire N__3274;
    wire N__3271;
    wire N__3268;
    wire N__3259;
    wire N__3258;
    wire N__3255;
    wire N__3254;
    wire N__3253;
    wire N__3250;
    wire N__3249;
    wire N__3246;
    wire N__3241;
    wire N__3236;
    wire N__3229;
    wire N__3226;
    wire N__3223;
    wire N__3220;
    wire N__3217;
    wire N__3214;
    wire N__3213;
    wire N__3212;
    wire N__3211;
    wire N__3208;
    wire N__3205;
    wire N__3200;
    wire N__3193;
    wire N__3192;
    wire N__3191;
    wire N__3188;
    wire N__3185;
    wire N__3182;
    wire N__3175;
    wire N__3172;
    wire N__3169;
    wire N__3166;
    wire N__3163;
    wire N__3160;
    wire N__3157;
    wire N__3154;
    wire N__3151;
    wire N__3148;
    wire N__3145;
    wire N__3142;
    wire N__3139;
    wire N__3136;
    wire N__3133;
    wire N__3130;
    wire N__3129;
    wire N__3126;
    wire N__3123;
    wire N__3120;
    wire N__3119;
    wire N__3116;
    wire N__3113;
    wire N__3110;
    wire N__3107;
    wire N__3104;
    wire N__3099;
    wire N__3094;
    wire N__3091;
    wire N__3088;
    wire N__3085;
    wire N__3082;
    wire N__3079;
    wire N__3076;
    wire N__3073;
    wire N__3070;
    wire N__3067;
    wire N__3064;
    wire N__3061;
    wire N__3058;
    wire N__3055;
    wire N__3052;
    wire N__3049;
    wire N__3046;
    wire N__3043;
    wire N__3040;
    wire N__3037;
    wire N__3034;
    wire N__3031;
    wire N__3028;
    wire N__3025;
    wire N__3022;
    wire N__3019;
    wire N__3016;
    wire N__3013;
    wire N__3010;
    wire N__3007;
    wire N__3004;
    wire N__3001;
    wire N__2998;
    wire N__2995;
    wire N__2992;
    wire N__2989;
    wire N__2986;
    wire N__2983;
    wire N__2980;
    wire N__2977;
    wire N__2974;
    wire N__2971;
    wire N__2970;
    wire N__2967;
    wire N__2964;
    wire N__2959;
    wire N__2956;
    wire N__2953;
    wire N__2950;
    wire N__2947;
    wire N__2944;
    wire N__2941;
    wire N__2938;
    wire N__2935;
    wire N__2932;
    wire N__2929;
    wire N__2926;
    wire N__2923;
    wire N__2920;
    wire N__2917;
    wire N__2914;
    wire N__2911;
    wire N__2908;
    wire N__2905;
    wire N__2902;
    wire N__2899;
    wire N__2896;
    wire N__2893;
    wire N__2892;
    wire N__2889;
    wire N__2886;
    wire N__2881;
    wire N__2878;
    wire N__2875;
    wire N__2872;
    wire N__2871;
    wire N__2868;
    wire N__2865;
    wire N__2860;
    wire N__2857;
    wire N__2854;
    wire N__2851;
    wire N__2848;
    wire N__2845;
    wire N__2842;
    wire N__2839;
    wire N__2838;
    wire N__2835;
    wire N__2832;
    wire N__2829;
    wire N__2826;
    wire N__2823;
    wire N__2818;
    wire N__2815;
    wire N__2812;
    wire N__2809;
    wire N__2806;
    wire N__2803;
    wire N__2800;
    wire N__2797;
    wire N__2794;
    wire N__2791;
    wire N__2788;
    wire N__2785;
    wire N__2782;
    wire N__2779;
    wire N__2776;
    wire N__2773;
    wire N__2770;
    wire N__2767;
    wire N__2764;
    wire N__2761;
    wire N__2758;
    wire N__2755;
    wire N__2752;
    wire N__2749;
    wire N__2746;
    wire VCCG0;
    wire clk_in_c;
    wire clk;
    wire GNDG0;
    wire uart_RXD;
    wire o_serial_data_c;
    wire bfn_6_11_0_;
    wire \Glue_Lab2.reset_count_cry_0 ;
    wire \Glue_Lab2.reset_count_cry_1 ;
    wire \Glue_Lab2.reset_count_cry_2 ;
    wire \Glue_Lab2.reset_count_cry_3 ;
    wire \Glue_Lab2.reset_count_cry_1_THRU_CO ;
    wire \Glue_Lab2.reset_countZ0Z_2 ;
    wire \buart.Z_tx.shifterZ0Z_1 ;
    wire \buart.Z_tx.shifterZ0Z_0 ;
    wire \buart.Z_tx.shifterZ0Z_2 ;
    wire \buart.Z_tx.shifterZ0Z_3 ;
    wire \buart.Z_tx.shifterZ0Z_4 ;
    wire \buart.Z_tx.shifterZ0Z_5 ;
    wire \buart.Z_tx.shifterZ0Z_7 ;
    wire \buart.Z_tx.shifterZ0Z_6 ;
    wire \Glue_Lab2.reset_count_cry_2_THRU_CO ;
    wire \Glue_Lab2.reset_countZ0Z_3 ;
    wire \Glue_Lab2.reset_count_cry_0_THRU_CO ;
    wire \Glue_Lab2.reset_countZ0Z_1 ;
    wire \buart.Z_rx.Z_baudgen.counter_0_1_5_cascade_ ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_ac0_7 ;
    wire \buart.Z_rx.ser_clk_2_cascade_ ;
    wire \Glue_Lab2.reset_countZ0Z_0 ;
    wire \buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_4 ;
    wire \Lab_UT.sDelay.delayRegZ0Z_0 ;
    wire Gl_tx_data_0;
    wire \Lab_UT.S_m_bmZ0Z_3_cascade_ ;
    wire led_c_3;
    wire led_c_3_cascade_;
    wire Gl_tx_data_3;
    wire \Lab_UT.S_m_bm_N_3LZ0Z3 ;
    wire \Lab_UT.g0_0_a3_0Z0Z_0_cascade_ ;
    wire Lab_UT_C_out41_1_cascade_;
    wire Gl_tx_data_5;
    wire \Lab_UT.N_6_0 ;
    wire \Lab_UT.g0_0_a3Z0Z_0_cascade_ ;
    wire \Lab_UT.g0_1Z0Z_0 ;
    wire \Lab_UT.N_6 ;
    wire \Lab_UT.S_0_s_axbZ0Z3_cascade_ ;
    wire \Lab_UT.S_m_amZ0Z_3 ;
    wire \Lab_UT.g1_0_0 ;
    wire \Lab_UT.S_m_bm_N_6LZ0Z10 ;
    wire \Glue_Lab2.g0_9_0_cascade_ ;
    wire \Glue_Lab2.reset_counte_0_1 ;
    wire \Glue_Lab2.g0_7_0 ;
    wire \buart.Z_rx.bitcountlde_0_cascade_ ;
    wire CONSTANT_ONE_NET;
    wire \buart.Z_rx.N_29_0_i_cascade_ ;
    wire \buart.Z_rx.bitcount_lm_0 ;
    wire \Glue_Lab2.de0.g0_5_0 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_0 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_1 ;
    wire \Glue_Lab2.de0.g0_5_2_cascade_ ;
    wire \Glue_Lab2.g0_9_2_cascade_ ;
    wire \Glue_Lab2.g0_7_2 ;
    wire \Glue_Lab2.reset_counte_0_3 ;
    wire \buart.Z_rx.bitcount_RNIMK771_0Z0Z_4_cascade_ ;
    wire bu_rx_data_rdy_cascade_;
    wire \Glue_Lab2.i_rst_char_detected ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_4 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_5 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_3 ;
    wire \buart.Z_rx.un1_sample_0 ;
    wire \buart.Z_rx.ser_clk_2_0_cascade_ ;
    wire \Glue_Lab2.de0.un2_de_hexplus_3_xZ0Z0_cascade_ ;
    wire \Glue_Lab2.de0.un2_de_hexplus_3_cascade_ ;
    wire \Glue_Lab2.is_hexplus_cascade_ ;
    wire Gl_tx_data_4;
    wire \buart.Z_rx.ser_clk_2 ;
    wire \buart.Z_rx.ser_clk_2_0 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_2 ;
    wire \Glue_Lab2.gl_fsm.N_14_cascade_ ;
    wire Glue_Lab2_gl_fsm_state_0;
    wire \Lab_UT.C_out41_0 ;
    wire led_c_0_4_cascade_;
    wire Gl_tx_data_6;
    wire \Lab_UT.S_m_bm_N_2LZ0Z1 ;
    wire led_c_0;
    wire \Lab_UT.S_1_ac0_1_0Z0Z_0 ;
    wire \Lab_UT.S_1_axbZ0Z1_cascade_ ;
    wire \Lab_UT.g1Z0Z_0 ;
    wire \Lab_UT.S_0_s_c2_0_cascade_ ;
    wire \Lab_UT.S_0_s_ac0_5_0_1 ;
    wire \Lab_UT.gZ0Z1 ;
    wire Glue_Lab2_Gl_r2_fast_0;
    wire Glue_Lab2_Gl_r1_fast_0;
    wire \Lab_UT.S_m_bm_N_5LZ0Z7 ;
    wire Gl_r1_2_rep1;
    wire Gl_r2_2_rep1;
    wire \Lab_UT.g0_4Z0Z_0 ;
    wire \Glue_Lab2.Gl_r17_0_i ;
    wire \Lab_UT.g0_1_0_0 ;
    wire \Glue_Lab2.Gl_r27_0_i ;
    wire \Lab_UT.g0_4_0_0 ;
    wire \Lab_UT.S_0_s_c2_1_cascade_ ;
    wire \Lab_UT.S_0_s_ac0_5_0_2 ;
    wire Lab_UT_g1_1;
    wire bfn_9_9_0_;
    wire \buart.Z_rx.bitcount_cry_0 ;
    wire \buart.Z_rx.bitcount_cry_1 ;
    wire \buart.Z_rx.bitcount_cry_2 ;
    wire \buart.Z_rx.bitcount_cry_3 ;
    wire \buart.Z_rx.bitcount_lm_4 ;
    wire \buart.Z_rx.bitcount_cry_0_THRU_CO ;
    wire \buart.Z_rx.bitcount_cry_2_THRU_CO ;
    wire \buart.Z_rx.bitcount_lm_3_cascade_ ;
    wire buart__rx_bitcount_4;
    wire buart__rx_bitcount_3;
    wire \buart.Z_rx.bitcount_RNIMK771Z0Z_4_cascade_ ;
    wire \buart.Z_rx.idle ;
    wire \buart.Z_rx.idle_cascade_ ;
    wire \buart.Z_rx.hhZ0Z_0 ;
    wire \buart.Z_rx.startbit_cascade_ ;
    wire \buart.Z_rx.bitcount_lm_1 ;
    wire buart__rx_bitcount_1;
    wire \buart.Z_rx.bitcount_cry_1_THRU_CO ;
    wire \buart.Z_rx.N_29_0_i ;
    wire \buart.Z_rx.bitcountlde_0 ;
    wire \buart.Z_rx.bitcount_lm_2_cascade_ ;
    wire \buart.Z_rx.startbit ;
    wire buart__rx_bitcount_2;
    wire \Glue_Lab2.g0_8_2 ;
    wire \Glue_Lab2.de0.un2_de_hexplusZ0Z_2 ;
    wire \Glue_Lab2.de0.un1_charDataZ0 ;
    wire buart__rx_shifter_fast_5;
    wire \buart.Z_rx.hhZ0Z_1 ;
    wire \Glue_Lab2.g0_8_0 ;
    wire \Glue_Lab2.de0.de_escZ0Z_3 ;
    wire \Glue_Lab2.gl_fsm.enOp_0_a2_1 ;
    wire \Glue_Lab2.gl_fsm.enOp_0_a2Z0Z_4 ;
    wire bu_rx_data_rdy;
    wire \Glue_Lab2.Gl_r1_2_1_cascade_ ;
    wire \Glue_Lab2.Gl_r1_2_2_cascade_ ;
    wire \Lab_UT.g0Z0Z_1 ;
    wire \Glue_Lab2.enOp ;
    wire Gl_tx_data_2;
    wire Glue_Lab2_gl_fsm_state_1;
    wire \Glue_Lab2.gl_fsm.enOp_0_a2_2 ;
    wire \Glue_Lab2.Gl_subtract_1_cascade_ ;
    wire \Lab_UT.S_0_s_axbZ0Z3 ;
    wire \Lab_UT.S_0_s_cZ0Z2 ;
    wire \Lab_UT.S_m_amZ0Z_2_cascade_ ;
    wire led_c_2;
    wire Gl_r1_0;
    wire Gl_r2_1;
    wire Gl_r2_0;
    wire Gl_r1_1;
    wire \Lab_UT.S_m_amZ0Z_1 ;
    wire \Lab_UT.S_m_bmZ0Z_1_cascade_ ;
    wire led_c_1;
    wire led_c_1_cascade_;
    wire Gl_tx_data_1;
    wire Gl_r2_fast_2;
    wire Gl_r1_fast_2;
    wire \Lab_UT.S_m_bm_1Z0Z_2 ;
    wire \Lab_UT.S_m_bmZ0Z_2 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_c5_cascade_ ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_c5 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_4 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_5 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_6 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_1 ;
    wire \buart.Z_tx.Z_baudgen.ser_clk_sx_cascade_ ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_0 ;
    wire \buart.Z_tx.Z_baudgen.counter_RNIES38_0Z0Z_4 ;
    wire \buart.Z_tx.Z_baudgen.un1_bitcount_c2_1 ;
    wire \buart.Z_tx.bitcount_RNIBADLZ0Z_1_cascade_ ;
    wire \buart.Z_tx.counter_RNIVE1P1_4_cascade_ ;
    wire \buart.Z_tx.un1_bitcount_c2 ;
    wire \buart.Z_tx.uart_busy_0_0 ;
    wire \buart.Z_tx.uart_busy_0_0_cascade_ ;
    wire \buart.Z_tx.bitcountZ0Z_2 ;
    wire \buart.Z_tx.un1_bitcount_c3_cascade_ ;
    wire \buart.Z_tx.bitcountZ0Z_3 ;
    wire \buart.Z_tx.un1_uart_wr_i_0_i_sx ;
    wire \Glue_Lab2.is_hexplus ;
    wire \buart.Z_tx.un1_bitcount_c1_cascade_ ;
    wire \buart.Z_tx.bitcountZ0Z_1 ;
    wire \buart.Z_tx.counter_RNIVE1P1_4 ;
    wire \buart.Z_tx.bitcountZ0Z_0 ;
    wire \Glue_Lab2.de0.de_escZ0Z_4 ;
    wire \Glue_Lab2.de0.g0_5_1_cascade_ ;
    wire \Glue_Lab2.g0_9_1_cascade_ ;
    wire \Glue_Lab2.g0_7_1 ;
    wire \Glue_Lab2.reset_counte_0_2 ;
    wire bu_rx_data_4;
    wire buart__rx_bitcount_0;
    wire \Glue_Lab2.de0.g0Z0Z_5_cascade_ ;
    wire bu_rx_data_0;
    wire \Glue_Lab2.reset_countZ0Z_4 ;
    wire \Glue_Lab2.g0_9_cascade_ ;
    wire \Glue_Lab2.g0_7 ;
    wire \Glue_Lab2.reset_counte_0_0 ;
    wire bu_rx_data_2;
    wire bu_rx_data_6;
    wire buart__rx_shifter_fast_4;
    wire \buart.Z_rx.sample ;
    wire Glue_Lab2_Gl_Op_0;
    wire Glue_Lab2_Gl_Op_3;
    wire Glue_Lab2_Gl_Op_1;
    wire Glue_Lab2_Gl_Op_5;
    wire \Glue_Lab2.g0_0_1_0_cascade_ ;
    wire Glue_Lab2_Gl_Op_2;
    wire \Glue_Lab2.Gl_subtract_0 ;
    wire Gl_r1_2;
    wire Gl_r2_2;
    wire Gl_r1_3;
    wire \Lab_UT.S_1_c3_d ;
    wire \Lab_UT.S_1_c3_cZ0_cascade_ ;
    wire Gl_r2_3;
    wire \Lab_UT.S_0_s_ac0_5_0Z0Z_0 ;
    wire \Lab_UT.S_0_s_ac0_5_dZ0 ;
    wire \Lab_UT.C_out41_cascade_ ;
    wire Gl_subtract;
    wire led_c_4;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_2 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_c2 ;
    wire \buart.Z_tx.ser_clk ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_3 ;
    wire Gl_tx_data_rdy;
    wire \buart.Z_tx.shifterZ0Z_8 ;
    wire \buart.Z_tx.un1_uart_wr_i_0_i ;
    wire \Glue_Lab2.g0_8 ;
    wire bu_rx_data_7;
    wire bu_rx_data_3;
    wire bu_rx_data_5;
    wire bu_rx_data_1;
    wire \Glue_Lab2.g0_8_1 ;
    wire \Lab_UT.sDelay.delayRegZ0Z_1 ;
    wire \Lab_UT.sDelay.delayRegZ0Z_2 ;
    wire \Lab_UT.sDelay.delayRegZ0Z_3 ;
    wire Gl_rst;
    wire L2_adder_rdy;
    wire clk_g;
    wire _gnd_net_;

    defparam ice_pll_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam ice_pll_inst.TEST_MODE=1'b0;
    defparam ice_pll_inst.SHIFTREG_DIV_MODE=2'b00;
    defparam ice_pll_inst.PLLOUT_SELECT="GENCLK";
    defparam ice_pll_inst.FILTER_RANGE=3'b001;
    defparam ice_pll_inst.FEEDBACK_PATH="SIMPLE";
    defparam ice_pll_inst.FDA_RELATIVE=4'b0000;
    defparam ice_pll_inst.FDA_FEEDBACK=4'b0000;
    defparam ice_pll_inst.ENABLE_ICEGATE=1'b0;
    defparam ice_pll_inst.DIVR=4'b0000;
    defparam ice_pll_inst.DIVQ=3'b100;
    defparam ice_pll_inst.DIVF=7'b0111111;
    defparam ice_pll_inst.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE ice_pll_inst (
            .EXTFEEDBACK(),
            .LATCHINPUTVALUE(),
            .SCLK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(clk),
            .REFERENCECLK(N__2806),
            .RESETB(N__3133),
            .BYPASS(GNDG0),
            .SDI(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    IO_PAD led_obuf_0_iopad (
            .OE(N__7037),
            .DIN(N__7036),
            .DOUT(N__7035),
            .PACKAGEPIN(led[0]));
    defparam led_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_0_preio (
            .PADOEN(N__7037),
            .PADOUT(N__7036),
            .PADIN(N__7035),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3469),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD test1_obuf_iopad (
            .OE(N__7028),
            .DIN(N__7027),
            .DOUT(N__7026),
            .PACKAGEPIN(test1));
    defparam test1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam test1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO test1_obuf_preio (
            .PADOEN(N__7028),
            .PADOUT(N__7027),
            .PADIN(N__7026),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD \Z_rcxd.Z_io_iopad  (
            .OE(N__7019),
            .DIN(N__7018),
            .DOUT(N__7017),
            .PACKAGEPIN(from_pc));
    defparam \Z_rcxd.Z_io_preio .PIN_TYPE=6'b000000;
    PRE_IO \Z_rcxd.Z_io_preio  (
            .PADOEN(N__7019),
            .PADOUT(N__7018),
            .PADIN(N__7017),
            .CLOCKENABLE(),
            .DOUT1(GNDG0),
            .OUTPUTENABLE(),
            .DIN0(uart_RXD),
            .DOUT0(GNDG0),
            .INPUTCLK(N__6162),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD sd_obuf_iopad (
            .OE(N__7010),
            .DIN(N__7009),
            .DOUT(N__7008),
            .PACKAGEPIN(sd));
    defparam sd_obuf_preio.NEG_TRIGGER=1'b0;
    defparam sd_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO sd_obuf_preio (
            .PADOEN(N__7010),
            .PADOUT(N__7009),
            .PADIN(N__7008),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD clk_in_ibuf_iopad (
            .OE(N__7001),
            .DIN(N__7000),
            .DOUT(N__6999),
            .PACKAGEPIN(clk_in));
    defparam clk_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam clk_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_in_ibuf_preio (
            .PADOEN(N__7001),
            .PADOUT(N__7000),
            .PADIN(N__6999),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(clk_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_2_iopad (
            .OE(N__6992),
            .DIN(N__6991),
            .DOUT(N__6990),
            .PACKAGEPIN(led[2]));
    defparam led_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_2_preio (
            .PADOEN(N__6992),
            .PADOUT(N__6991),
            .PADIN(N__6990),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4621),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_4_iopad (
            .OE(N__6983),
            .DIN(N__6982),
            .DOUT(N__6981),
            .PACKAGEPIN(led[4]));
    defparam led_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_4_preio (
            .PADOEN(N__6983),
            .PADOUT(N__6982),
            .PADIN(N__6981),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5542),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD test3_obuf_iopad (
            .OE(N__6974),
            .DIN(N__6973),
            .DOUT(N__6972),
            .PACKAGEPIN(test3));
    defparam test3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam test3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO test3_obuf_preio (
            .PADOEN(N__6974),
            .PADOUT(N__6973),
            .PADIN(N__6972),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD to_ir_obuf_iopad (
            .OE(N__6965),
            .DIN(N__6964),
            .DOUT(N__6963),
            .PACKAGEPIN(to_ir));
    defparam to_ir_obuf_preio.NEG_TRIGGER=1'b0;
    defparam to_ir_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO to_ir_obuf_preio (
            .PADOEN(N__6965),
            .PADOUT(N__6964),
            .PADIN(N__6963),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_1_iopad (
            .OE(N__6956),
            .DIN(N__6955),
            .DOUT(N__6954),
            .PACKAGEPIN(led[1]));
    defparam led_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_1_preio (
            .PADOEN(N__6956),
            .PADOUT(N__6955),
            .PADIN(N__6954),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4342),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_3_iopad (
            .OE(N__6947),
            .DIN(N__6946),
            .DOUT(N__6945),
            .PACKAGEPIN(led[3]));
    defparam led_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_3_preio (
            .PADOEN(N__6947),
            .PADOUT(N__6946),
            .PADIN(N__6945),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3034),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_serial_data_obuf_iopad (
            .OE(N__6938),
            .DIN(N__6937),
            .DOUT(N__6936),
            .PACKAGEPIN(o_serial_data));
    defparam o_serial_data_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_serial_data_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_serial_data_obuf_preio (
            .PADOEN(N__6938),
            .PADOUT(N__6937),
            .PADIN(N__6936),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2761),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD test2_obuf_iopad (
            .OE(N__6929),
            .DIN(N__6928),
            .DOUT(N__6927),
            .PACKAGEPIN(test2));
    defparam test2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam test2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO test2_obuf_preio (
            .PADOEN(N__6929),
            .PADOUT(N__6928),
            .PADIN(N__6927),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__1620 (
            .O(N__6910),
            .I(N__6900));
    InMux I__1619 (
            .O(N__6909),
            .I(N__6900));
    InMux I__1618 (
            .O(N__6908),
            .I(N__6891));
    InMux I__1617 (
            .O(N__6907),
            .I(N__6891));
    InMux I__1616 (
            .O(N__6906),
            .I(N__6891));
    InMux I__1615 (
            .O(N__6905),
            .I(N__6891));
    LocalMux I__1614 (
            .O(N__6900),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ));
    LocalMux I__1613 (
            .O(N__6891),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ));
    CascadeMux I__1612 (
            .O(N__6886),
            .I(N__6882));
    CascadeMux I__1611 (
            .O(N__6885),
            .I(N__6878));
    InMux I__1610 (
            .O(N__6882),
            .I(N__6872));
    InMux I__1609 (
            .O(N__6881),
            .I(N__6872));
    InMux I__1608 (
            .O(N__6878),
            .I(N__6867));
    InMux I__1607 (
            .O(N__6877),
            .I(N__6867));
    LocalMux I__1606 (
            .O(N__6872),
            .I(N__6864));
    LocalMux I__1605 (
            .O(N__6867),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_c2 ));
    Odrv4 I__1604 (
            .O(N__6864),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_c2 ));
    InMux I__1603 (
            .O(N__6859),
            .I(N__6850));
    InMux I__1602 (
            .O(N__6858),
            .I(N__6850));
    InMux I__1601 (
            .O(N__6857),
            .I(N__6845));
    InMux I__1600 (
            .O(N__6856),
            .I(N__6840));
    InMux I__1599 (
            .O(N__6855),
            .I(N__6840));
    LocalMux I__1598 (
            .O(N__6850),
            .I(N__6837));
    InMux I__1597 (
            .O(N__6849),
            .I(N__6832));
    InMux I__1596 (
            .O(N__6848),
            .I(N__6832));
    LocalMux I__1595 (
            .O(N__6845),
            .I(\buart.Z_tx.ser_clk ));
    LocalMux I__1594 (
            .O(N__6840),
            .I(\buart.Z_tx.ser_clk ));
    Odrv4 I__1593 (
            .O(N__6837),
            .I(\buart.Z_tx.ser_clk ));
    LocalMux I__1592 (
            .O(N__6832),
            .I(\buart.Z_tx.ser_clk ));
    CascadeMux I__1591 (
            .O(N__6823),
            .I(N__6817));
    CascadeMux I__1590 (
            .O(N__6822),
            .I(N__6814));
    InMux I__1589 (
            .O(N__6821),
            .I(N__6810));
    InMux I__1588 (
            .O(N__6820),
            .I(N__6801));
    InMux I__1587 (
            .O(N__6817),
            .I(N__6801));
    InMux I__1586 (
            .O(N__6814),
            .I(N__6801));
    InMux I__1585 (
            .O(N__6813),
            .I(N__6801));
    LocalMux I__1584 (
            .O(N__6810),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ));
    LocalMux I__1583 (
            .O(N__6801),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ));
    InMux I__1582 (
            .O(N__6796),
            .I(N__6782));
    InMux I__1581 (
            .O(N__6795),
            .I(N__6765));
    InMux I__1580 (
            .O(N__6794),
            .I(N__6765));
    InMux I__1579 (
            .O(N__6793),
            .I(N__6765));
    InMux I__1578 (
            .O(N__6792),
            .I(N__6765));
    InMux I__1577 (
            .O(N__6791),
            .I(N__6765));
    InMux I__1576 (
            .O(N__6790),
            .I(N__6765));
    InMux I__1575 (
            .O(N__6789),
            .I(N__6765));
    InMux I__1574 (
            .O(N__6788),
            .I(N__6765));
    InMux I__1573 (
            .O(N__6787),
            .I(N__6754));
    InMux I__1572 (
            .O(N__6786),
            .I(N__6754));
    InMux I__1571 (
            .O(N__6785),
            .I(N__6754));
    LocalMux I__1570 (
            .O(N__6782),
            .I(N__6749));
    LocalMux I__1569 (
            .O(N__6765),
            .I(N__6749));
    InMux I__1568 (
            .O(N__6764),
            .I(N__6746));
    InMux I__1567 (
            .O(N__6763),
            .I(N__6739));
    InMux I__1566 (
            .O(N__6762),
            .I(N__6739));
    InMux I__1565 (
            .O(N__6761),
            .I(N__6739));
    LocalMux I__1564 (
            .O(N__6754),
            .I(N__6736));
    Odrv12 I__1563 (
            .O(N__6749),
            .I(Gl_tx_data_rdy));
    LocalMux I__1562 (
            .O(N__6746),
            .I(Gl_tx_data_rdy));
    LocalMux I__1561 (
            .O(N__6739),
            .I(Gl_tx_data_rdy));
    Odrv4 I__1560 (
            .O(N__6736),
            .I(Gl_tx_data_rdy));
    InMux I__1559 (
            .O(N__6727),
            .I(N__6724));
    LocalMux I__1558 (
            .O(N__6724),
            .I(N__6721));
    Span4Mux_h I__1557 (
            .O(N__6721),
            .I(N__6718));
    Odrv4 I__1556 (
            .O(N__6718),
            .I(\buart.Z_tx.shifterZ0Z_8 ));
    CEMux I__1555 (
            .O(N__6715),
            .I(N__6712));
    LocalMux I__1554 (
            .O(N__6712),
            .I(N__6708));
    CEMux I__1553 (
            .O(N__6711),
            .I(N__6705));
    Span4Mux_h I__1552 (
            .O(N__6708),
            .I(N__6702));
    LocalMux I__1551 (
            .O(N__6705),
            .I(N__6698));
    Span4Mux_s1_h I__1550 (
            .O(N__6702),
            .I(N__6695));
    CEMux I__1549 (
            .O(N__6701),
            .I(N__6692));
    Odrv12 I__1548 (
            .O(N__6698),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i ));
    Odrv4 I__1547 (
            .O(N__6695),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i ));
    LocalMux I__1546 (
            .O(N__6692),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i ));
    InMux I__1545 (
            .O(N__6685),
            .I(N__6682));
    LocalMux I__1544 (
            .O(N__6682),
            .I(\Glue_Lab2.g0_8 ));
    InMux I__1543 (
            .O(N__6679),
            .I(N__6676));
    LocalMux I__1542 (
            .O(N__6676),
            .I(N__6669));
    InMux I__1541 (
            .O(N__6675),
            .I(N__6666));
    InMux I__1540 (
            .O(N__6674),
            .I(N__6663));
    CascadeMux I__1539 (
            .O(N__6673),
            .I(N__6656));
    CascadeMux I__1538 (
            .O(N__6672),
            .I(N__6653));
    Span4Mux_s2_h I__1537 (
            .O(N__6669),
            .I(N__6650));
    LocalMux I__1536 (
            .O(N__6666),
            .I(N__6647));
    LocalMux I__1535 (
            .O(N__6663),
            .I(N__6644));
    InMux I__1534 (
            .O(N__6662),
            .I(N__6639));
    InMux I__1533 (
            .O(N__6661),
            .I(N__6639));
    InMux I__1532 (
            .O(N__6660),
            .I(N__6630));
    InMux I__1531 (
            .O(N__6659),
            .I(N__6630));
    InMux I__1530 (
            .O(N__6656),
            .I(N__6630));
    InMux I__1529 (
            .O(N__6653),
            .I(N__6630));
    Odrv4 I__1528 (
            .O(N__6650),
            .I(bu_rx_data_7));
    Odrv12 I__1527 (
            .O(N__6647),
            .I(bu_rx_data_7));
    Odrv4 I__1526 (
            .O(N__6644),
            .I(bu_rx_data_7));
    LocalMux I__1525 (
            .O(N__6639),
            .I(bu_rx_data_7));
    LocalMux I__1524 (
            .O(N__6630),
            .I(bu_rx_data_7));
    InMux I__1523 (
            .O(N__6619),
            .I(N__6616));
    LocalMux I__1522 (
            .O(N__6616),
            .I(N__6609));
    InMux I__1521 (
            .O(N__6615),
            .I(N__6606));
    InMux I__1520 (
            .O(N__6614),
            .I(N__6603));
    InMux I__1519 (
            .O(N__6613),
            .I(N__6600));
    InMux I__1518 (
            .O(N__6612),
            .I(N__6597));
    Span4Mux_s1_v I__1517 (
            .O(N__6609),
            .I(N__6590));
    LocalMux I__1516 (
            .O(N__6606),
            .I(N__6590));
    LocalMux I__1515 (
            .O(N__6603),
            .I(N__6587));
    LocalMux I__1514 (
            .O(N__6600),
            .I(N__6582));
    LocalMux I__1513 (
            .O(N__6597),
            .I(N__6582));
    InMux I__1512 (
            .O(N__6596),
            .I(N__6579));
    CascadeMux I__1511 (
            .O(N__6595),
            .I(N__6573));
    Span4Mux_v I__1510 (
            .O(N__6590),
            .I(N__6569));
    Span4Mux_h I__1509 (
            .O(N__6587),
            .I(N__6566));
    Span4Mux_s2_h I__1508 (
            .O(N__6582),
            .I(N__6563));
    LocalMux I__1507 (
            .O(N__6579),
            .I(N__6560));
    InMux I__1506 (
            .O(N__6578),
            .I(N__6555));
    InMux I__1505 (
            .O(N__6577),
            .I(N__6555));
    InMux I__1504 (
            .O(N__6576),
            .I(N__6548));
    InMux I__1503 (
            .O(N__6573),
            .I(N__6548));
    InMux I__1502 (
            .O(N__6572),
            .I(N__6548));
    Odrv4 I__1501 (
            .O(N__6569),
            .I(bu_rx_data_3));
    Odrv4 I__1500 (
            .O(N__6566),
            .I(bu_rx_data_3));
    Odrv4 I__1499 (
            .O(N__6563),
            .I(bu_rx_data_3));
    Odrv4 I__1498 (
            .O(N__6560),
            .I(bu_rx_data_3));
    LocalMux I__1497 (
            .O(N__6555),
            .I(bu_rx_data_3));
    LocalMux I__1496 (
            .O(N__6548),
            .I(bu_rx_data_3));
    CascadeMux I__1495 (
            .O(N__6535),
            .I(N__6531));
    CascadeMux I__1494 (
            .O(N__6534),
            .I(N__6525));
    InMux I__1493 (
            .O(N__6531),
            .I(N__6520));
    InMux I__1492 (
            .O(N__6530),
            .I(N__6520));
    CascadeMux I__1491 (
            .O(N__6529),
            .I(N__6516));
    CascadeMux I__1490 (
            .O(N__6528),
            .I(N__6513));
    InMux I__1489 (
            .O(N__6525),
            .I(N__6510));
    LocalMux I__1488 (
            .O(N__6520),
            .I(N__6507));
    InMux I__1487 (
            .O(N__6519),
            .I(N__6502));
    InMux I__1486 (
            .O(N__6516),
            .I(N__6499));
    InMux I__1485 (
            .O(N__6513),
            .I(N__6496));
    LocalMux I__1484 (
            .O(N__6510),
            .I(N__6491));
    Span4Mux_v I__1483 (
            .O(N__6507),
            .I(N__6491));
    InMux I__1482 (
            .O(N__6506),
            .I(N__6486));
    InMux I__1481 (
            .O(N__6505),
            .I(N__6486));
    LocalMux I__1480 (
            .O(N__6502),
            .I(bu_rx_data_5));
    LocalMux I__1479 (
            .O(N__6499),
            .I(bu_rx_data_5));
    LocalMux I__1478 (
            .O(N__6496),
            .I(bu_rx_data_5));
    Odrv4 I__1477 (
            .O(N__6491),
            .I(bu_rx_data_5));
    LocalMux I__1476 (
            .O(N__6486),
            .I(bu_rx_data_5));
    InMux I__1475 (
            .O(N__6475),
            .I(N__6466));
    InMux I__1474 (
            .O(N__6474),
            .I(N__6463));
    InMux I__1473 (
            .O(N__6473),
            .I(N__6457));
    InMux I__1472 (
            .O(N__6472),
            .I(N__6454));
    CascadeMux I__1471 (
            .O(N__6471),
            .I(N__6451));
    InMux I__1470 (
            .O(N__6470),
            .I(N__6447));
    CascadeMux I__1469 (
            .O(N__6469),
            .I(N__6443));
    LocalMux I__1468 (
            .O(N__6466),
            .I(N__6438));
    LocalMux I__1467 (
            .O(N__6463),
            .I(N__6438));
    InMux I__1466 (
            .O(N__6462),
            .I(N__6431));
    InMux I__1465 (
            .O(N__6461),
            .I(N__6431));
    InMux I__1464 (
            .O(N__6460),
            .I(N__6431));
    LocalMux I__1463 (
            .O(N__6457),
            .I(N__6428));
    LocalMux I__1462 (
            .O(N__6454),
            .I(N__6425));
    InMux I__1461 (
            .O(N__6451),
            .I(N__6422));
    InMux I__1460 (
            .O(N__6450),
            .I(N__6419));
    LocalMux I__1459 (
            .O(N__6447),
            .I(N__6416));
    InMux I__1458 (
            .O(N__6446),
            .I(N__6413));
    InMux I__1457 (
            .O(N__6443),
            .I(N__6410));
    Span4Mux_v I__1456 (
            .O(N__6438),
            .I(N__6399));
    LocalMux I__1455 (
            .O(N__6431),
            .I(N__6399));
    Span4Mux_s0_h I__1454 (
            .O(N__6428),
            .I(N__6399));
    Span4Mux_v I__1453 (
            .O(N__6425),
            .I(N__6399));
    LocalMux I__1452 (
            .O(N__6422),
            .I(N__6399));
    LocalMux I__1451 (
            .O(N__6419),
            .I(bu_rx_data_1));
    Odrv12 I__1450 (
            .O(N__6416),
            .I(bu_rx_data_1));
    LocalMux I__1449 (
            .O(N__6413),
            .I(bu_rx_data_1));
    LocalMux I__1448 (
            .O(N__6410),
            .I(bu_rx_data_1));
    Odrv4 I__1447 (
            .O(N__6399),
            .I(bu_rx_data_1));
    InMux I__1446 (
            .O(N__6388),
            .I(N__6385));
    LocalMux I__1445 (
            .O(N__6385),
            .I(\Glue_Lab2.g0_8_1 ));
    InMux I__1444 (
            .O(N__6382),
            .I(N__6379));
    LocalMux I__1443 (
            .O(N__6379),
            .I(N__6376));
    Odrv12 I__1442 (
            .O(N__6376),
            .I(\Lab_UT.sDelay.delayRegZ0Z_1 ));
    InMux I__1441 (
            .O(N__6373),
            .I(N__6370));
    LocalMux I__1440 (
            .O(N__6370),
            .I(\Lab_UT.sDelay.delayRegZ0Z_2 ));
    InMux I__1439 (
            .O(N__6367),
            .I(N__6364));
    LocalMux I__1438 (
            .O(N__6364),
            .I(\Lab_UT.sDelay.delayRegZ0Z_3 ));
    CascadeMux I__1437 (
            .O(N__6361),
            .I(N__6349));
    CascadeMux I__1436 (
            .O(N__6360),
            .I(N__6345));
    CascadeMux I__1435 (
            .O(N__6359),
            .I(N__6340));
    InMux I__1434 (
            .O(N__6358),
            .I(N__6333));
    InMux I__1433 (
            .O(N__6357),
            .I(N__6324));
    InMux I__1432 (
            .O(N__6356),
            .I(N__6324));
    InMux I__1431 (
            .O(N__6355),
            .I(N__6324));
    InMux I__1430 (
            .O(N__6354),
            .I(N__6324));
    InMux I__1429 (
            .O(N__6353),
            .I(N__6319));
    InMux I__1428 (
            .O(N__6352),
            .I(N__6319));
    InMux I__1427 (
            .O(N__6349),
            .I(N__6314));
    InMux I__1426 (
            .O(N__6348),
            .I(N__6314));
    InMux I__1425 (
            .O(N__6345),
            .I(N__6301));
    InMux I__1424 (
            .O(N__6344),
            .I(N__6301));
    InMux I__1423 (
            .O(N__6343),
            .I(N__6292));
    InMux I__1422 (
            .O(N__6340),
            .I(N__6292));
    InMux I__1421 (
            .O(N__6339),
            .I(N__6292));
    InMux I__1420 (
            .O(N__6338),
            .I(N__6292));
    InMux I__1419 (
            .O(N__6337),
            .I(N__6286));
    InMux I__1418 (
            .O(N__6336),
            .I(N__6286));
    LocalMux I__1417 (
            .O(N__6333),
            .I(N__6277));
    LocalMux I__1416 (
            .O(N__6324),
            .I(N__6277));
    LocalMux I__1415 (
            .O(N__6319),
            .I(N__6277));
    LocalMux I__1414 (
            .O(N__6314),
            .I(N__6277));
    InMux I__1413 (
            .O(N__6313),
            .I(N__6266));
    InMux I__1412 (
            .O(N__6312),
            .I(N__6266));
    InMux I__1411 (
            .O(N__6311),
            .I(N__6266));
    InMux I__1410 (
            .O(N__6310),
            .I(N__6266));
    InMux I__1409 (
            .O(N__6309),
            .I(N__6266));
    InMux I__1408 (
            .O(N__6308),
            .I(N__6259));
    InMux I__1407 (
            .O(N__6307),
            .I(N__6259));
    InMux I__1406 (
            .O(N__6306),
            .I(N__6259));
    LocalMux I__1405 (
            .O(N__6301),
            .I(N__6256));
    LocalMux I__1404 (
            .O(N__6292),
            .I(N__6253));
    InMux I__1403 (
            .O(N__6291),
            .I(N__6250));
    LocalMux I__1402 (
            .O(N__6286),
            .I(N__6239));
    Span4Mux_s3_v I__1401 (
            .O(N__6277),
            .I(N__6239));
    LocalMux I__1400 (
            .O(N__6266),
            .I(N__6239));
    LocalMux I__1399 (
            .O(N__6259),
            .I(N__6236));
    Span4Mux_s1_v I__1398 (
            .O(N__6256),
            .I(N__6229));
    Span4Mux_h I__1397 (
            .O(N__6253),
            .I(N__6229));
    LocalMux I__1396 (
            .O(N__6250),
            .I(N__6229));
    InMux I__1395 (
            .O(N__6249),
            .I(N__6226));
    InMux I__1394 (
            .O(N__6248),
            .I(N__6223));
    InMux I__1393 (
            .O(N__6247),
            .I(N__6218));
    InMux I__1392 (
            .O(N__6246),
            .I(N__6218));
    Span4Mux_h I__1391 (
            .O(N__6239),
            .I(N__6215));
    Odrv12 I__1390 (
            .O(N__6236),
            .I(Gl_rst));
    Odrv4 I__1389 (
            .O(N__6229),
            .I(Gl_rst));
    LocalMux I__1388 (
            .O(N__6226),
            .I(Gl_rst));
    LocalMux I__1387 (
            .O(N__6223),
            .I(Gl_rst));
    LocalMux I__1386 (
            .O(N__6218),
            .I(Gl_rst));
    Odrv4 I__1385 (
            .O(N__6215),
            .I(Gl_rst));
    InMux I__1384 (
            .O(N__6202),
            .I(N__6199));
    LocalMux I__1383 (
            .O(N__6199),
            .I(N__6196));
    Odrv4 I__1382 (
            .O(N__6196),
            .I(L2_adder_rdy));
    ClkMux I__1381 (
            .O(N__6193),
            .I(N__6097));
    ClkMux I__1380 (
            .O(N__6192),
            .I(N__6097));
    ClkMux I__1379 (
            .O(N__6191),
            .I(N__6097));
    ClkMux I__1378 (
            .O(N__6190),
            .I(N__6097));
    ClkMux I__1377 (
            .O(N__6189),
            .I(N__6097));
    ClkMux I__1376 (
            .O(N__6188),
            .I(N__6097));
    ClkMux I__1375 (
            .O(N__6187),
            .I(N__6097));
    ClkMux I__1374 (
            .O(N__6186),
            .I(N__6097));
    ClkMux I__1373 (
            .O(N__6185),
            .I(N__6097));
    ClkMux I__1372 (
            .O(N__6184),
            .I(N__6097));
    ClkMux I__1371 (
            .O(N__6183),
            .I(N__6097));
    ClkMux I__1370 (
            .O(N__6182),
            .I(N__6097));
    ClkMux I__1369 (
            .O(N__6181),
            .I(N__6097));
    ClkMux I__1368 (
            .O(N__6180),
            .I(N__6097));
    ClkMux I__1367 (
            .O(N__6179),
            .I(N__6097));
    ClkMux I__1366 (
            .O(N__6178),
            .I(N__6097));
    ClkMux I__1365 (
            .O(N__6177),
            .I(N__6097));
    ClkMux I__1364 (
            .O(N__6176),
            .I(N__6097));
    ClkMux I__1363 (
            .O(N__6175),
            .I(N__6097));
    ClkMux I__1362 (
            .O(N__6174),
            .I(N__6097));
    ClkMux I__1361 (
            .O(N__6173),
            .I(N__6097));
    ClkMux I__1360 (
            .O(N__6172),
            .I(N__6097));
    ClkMux I__1359 (
            .O(N__6171),
            .I(N__6097));
    ClkMux I__1358 (
            .O(N__6170),
            .I(N__6097));
    ClkMux I__1357 (
            .O(N__6169),
            .I(N__6097));
    ClkMux I__1356 (
            .O(N__6168),
            .I(N__6097));
    ClkMux I__1355 (
            .O(N__6167),
            .I(N__6097));
    ClkMux I__1354 (
            .O(N__6166),
            .I(N__6097));
    ClkMux I__1353 (
            .O(N__6165),
            .I(N__6097));
    ClkMux I__1352 (
            .O(N__6164),
            .I(N__6097));
    ClkMux I__1351 (
            .O(N__6163),
            .I(N__6097));
    ClkMux I__1350 (
            .O(N__6162),
            .I(N__6097));
    GlobalMux I__1349 (
            .O(N__6097),
            .I(N__6094));
    gio2CtrlBuf I__1348 (
            .O(N__6094),
            .I(clk_g));
    InMux I__1347 (
            .O(N__6091),
            .I(N__6087));
    InMux I__1346 (
            .O(N__6090),
            .I(N__6084));
    LocalMux I__1345 (
            .O(N__6087),
            .I(N__6081));
    LocalMux I__1344 (
            .O(N__6084),
            .I(N__6076));
    Span4Mux_v I__1343 (
            .O(N__6081),
            .I(N__6076));
    Odrv4 I__1342 (
            .O(N__6076),
            .I(buart__rx_shifter_fast_4));
    CEMux I__1341 (
            .O(N__6073),
            .I(N__6068));
    CEMux I__1340 (
            .O(N__6072),
            .I(N__6065));
    CEMux I__1339 (
            .O(N__6071),
            .I(N__6062));
    LocalMux I__1338 (
            .O(N__6068),
            .I(N__6059));
    LocalMux I__1337 (
            .O(N__6065),
            .I(N__6055));
    LocalMux I__1336 (
            .O(N__6062),
            .I(N__6052));
    Span4Mux_v I__1335 (
            .O(N__6059),
            .I(N__6049));
    CEMux I__1334 (
            .O(N__6058),
            .I(N__6046));
    Span4Mux_v I__1333 (
            .O(N__6055),
            .I(N__6041));
    Span4Mux_s1_h I__1332 (
            .O(N__6052),
            .I(N__6041));
    Span4Mux_s2_v I__1331 (
            .O(N__6049),
            .I(N__6036));
    LocalMux I__1330 (
            .O(N__6046),
            .I(N__6036));
    Odrv4 I__1329 (
            .O(N__6041),
            .I(\buart.Z_rx.sample ));
    Odrv4 I__1328 (
            .O(N__6036),
            .I(\buart.Z_rx.sample ));
    InMux I__1327 (
            .O(N__6031),
            .I(N__6026));
    InMux I__1326 (
            .O(N__6030),
            .I(N__6020));
    InMux I__1325 (
            .O(N__6029),
            .I(N__6020));
    LocalMux I__1324 (
            .O(N__6026),
            .I(N__6017));
    InMux I__1323 (
            .O(N__6025),
            .I(N__6014));
    LocalMux I__1322 (
            .O(N__6020),
            .I(Glue_Lab2_Gl_Op_0));
    Odrv12 I__1321 (
            .O(N__6017),
            .I(Glue_Lab2_Gl_Op_0));
    LocalMux I__1320 (
            .O(N__6014),
            .I(Glue_Lab2_Gl_Op_0));
    InMux I__1319 (
            .O(N__6007),
            .I(N__6002));
    InMux I__1318 (
            .O(N__6006),
            .I(N__5996));
    InMux I__1317 (
            .O(N__6005),
            .I(N__5996));
    LocalMux I__1316 (
            .O(N__6002),
            .I(N__5993));
    InMux I__1315 (
            .O(N__6001),
            .I(N__5990));
    LocalMux I__1314 (
            .O(N__5996),
            .I(Glue_Lab2_Gl_Op_3));
    Odrv4 I__1313 (
            .O(N__5993),
            .I(Glue_Lab2_Gl_Op_3));
    LocalMux I__1312 (
            .O(N__5990),
            .I(Glue_Lab2_Gl_Op_3));
    InMux I__1311 (
            .O(N__5983),
            .I(N__5978));
    CascadeMux I__1310 (
            .O(N__5982),
            .I(N__5974));
    InMux I__1309 (
            .O(N__5981),
            .I(N__5971));
    LocalMux I__1308 (
            .O(N__5978),
            .I(N__5968));
    InMux I__1307 (
            .O(N__5977),
            .I(N__5963));
    InMux I__1306 (
            .O(N__5974),
            .I(N__5963));
    LocalMux I__1305 (
            .O(N__5971),
            .I(N__5960));
    Odrv4 I__1304 (
            .O(N__5968),
            .I(Glue_Lab2_Gl_Op_1));
    LocalMux I__1303 (
            .O(N__5963),
            .I(Glue_Lab2_Gl_Op_1));
    Odrv4 I__1302 (
            .O(N__5960),
            .I(Glue_Lab2_Gl_Op_1));
    InMux I__1301 (
            .O(N__5953),
            .I(N__5947));
    InMux I__1300 (
            .O(N__5952),
            .I(N__5944));
    InMux I__1299 (
            .O(N__5951),
            .I(N__5941));
    InMux I__1298 (
            .O(N__5950),
            .I(N__5938));
    LocalMux I__1297 (
            .O(N__5947),
            .I(N__5935));
    LocalMux I__1296 (
            .O(N__5944),
            .I(N__5932));
    LocalMux I__1295 (
            .O(N__5941),
            .I(Glue_Lab2_Gl_Op_5));
    LocalMux I__1294 (
            .O(N__5938),
            .I(Glue_Lab2_Gl_Op_5));
    Odrv4 I__1293 (
            .O(N__5935),
            .I(Glue_Lab2_Gl_Op_5));
    Odrv4 I__1292 (
            .O(N__5932),
            .I(Glue_Lab2_Gl_Op_5));
    CascadeMux I__1291 (
            .O(N__5923),
            .I(\Glue_Lab2.g0_0_1_0_cascade_ ));
    InMux I__1290 (
            .O(N__5920),
            .I(N__5917));
    LocalMux I__1289 (
            .O(N__5917),
            .I(N__5911));
    InMux I__1288 (
            .O(N__5916),
            .I(N__5906));
    InMux I__1287 (
            .O(N__5915),
            .I(N__5906));
    InMux I__1286 (
            .O(N__5914),
            .I(N__5903));
    Odrv12 I__1285 (
            .O(N__5911),
            .I(Glue_Lab2_Gl_Op_2));
    LocalMux I__1284 (
            .O(N__5906),
            .I(Glue_Lab2_Gl_Op_2));
    LocalMux I__1283 (
            .O(N__5903),
            .I(Glue_Lab2_Gl_Op_2));
    InMux I__1282 (
            .O(N__5896),
            .I(N__5893));
    LocalMux I__1281 (
            .O(N__5893),
            .I(N__5890));
    Span4Mux_h I__1280 (
            .O(N__5890),
            .I(N__5887));
    Odrv4 I__1279 (
            .O(N__5887),
            .I(\Glue_Lab2.Gl_subtract_0 ));
    InMux I__1278 (
            .O(N__5884),
            .I(N__5877));
    InMux I__1277 (
            .O(N__5883),
            .I(N__5877));
    InMux I__1276 (
            .O(N__5882),
            .I(N__5874));
    LocalMux I__1275 (
            .O(N__5877),
            .I(N__5868));
    LocalMux I__1274 (
            .O(N__5874),
            .I(N__5865));
    InMux I__1273 (
            .O(N__5873),
            .I(N__5857));
    InMux I__1272 (
            .O(N__5872),
            .I(N__5854));
    InMux I__1271 (
            .O(N__5871),
            .I(N__5851));
    Span4Mux_h I__1270 (
            .O(N__5868),
            .I(N__5846));
    Span4Mux_h I__1269 (
            .O(N__5865),
            .I(N__5846));
    InMux I__1268 (
            .O(N__5864),
            .I(N__5841));
    InMux I__1267 (
            .O(N__5863),
            .I(N__5841));
    InMux I__1266 (
            .O(N__5862),
            .I(N__5836));
    InMux I__1265 (
            .O(N__5861),
            .I(N__5836));
    InMux I__1264 (
            .O(N__5860),
            .I(N__5833));
    LocalMux I__1263 (
            .O(N__5857),
            .I(N__5830));
    LocalMux I__1262 (
            .O(N__5854),
            .I(Gl_r1_2));
    LocalMux I__1261 (
            .O(N__5851),
            .I(Gl_r1_2));
    Odrv4 I__1260 (
            .O(N__5846),
            .I(Gl_r1_2));
    LocalMux I__1259 (
            .O(N__5841),
            .I(Gl_r1_2));
    LocalMux I__1258 (
            .O(N__5836),
            .I(Gl_r1_2));
    LocalMux I__1257 (
            .O(N__5833),
            .I(Gl_r1_2));
    Odrv4 I__1256 (
            .O(N__5830),
            .I(Gl_r1_2));
    InMux I__1255 (
            .O(N__5815),
            .I(N__5806));
    InMux I__1254 (
            .O(N__5814),
            .I(N__5806));
    InMux I__1253 (
            .O(N__5813),
            .I(N__5802));
    CascadeMux I__1252 (
            .O(N__5812),
            .I(N__5797));
    CascadeMux I__1251 (
            .O(N__5811),
            .I(N__5794));
    LocalMux I__1250 (
            .O(N__5806),
            .I(N__5791));
    InMux I__1249 (
            .O(N__5805),
            .I(N__5788));
    LocalMux I__1248 (
            .O(N__5802),
            .I(N__5785));
    CascadeMux I__1247 (
            .O(N__5801),
            .I(N__5781));
    InMux I__1246 (
            .O(N__5800),
            .I(N__5776));
    InMux I__1245 (
            .O(N__5797),
            .I(N__5773));
    InMux I__1244 (
            .O(N__5794),
            .I(N__5770));
    Span4Mux_h I__1243 (
            .O(N__5791),
            .I(N__5763));
    LocalMux I__1242 (
            .O(N__5788),
            .I(N__5763));
    Span4Mux_h I__1241 (
            .O(N__5785),
            .I(N__5763));
    InMux I__1240 (
            .O(N__5784),
            .I(N__5760));
    InMux I__1239 (
            .O(N__5781),
            .I(N__5757));
    InMux I__1238 (
            .O(N__5780),
            .I(N__5752));
    InMux I__1237 (
            .O(N__5779),
            .I(N__5752));
    LocalMux I__1236 (
            .O(N__5776),
            .I(N__5749));
    LocalMux I__1235 (
            .O(N__5773),
            .I(Gl_r2_2));
    LocalMux I__1234 (
            .O(N__5770),
            .I(Gl_r2_2));
    Odrv4 I__1233 (
            .O(N__5763),
            .I(Gl_r2_2));
    LocalMux I__1232 (
            .O(N__5760),
            .I(Gl_r2_2));
    LocalMux I__1231 (
            .O(N__5757),
            .I(Gl_r2_2));
    LocalMux I__1230 (
            .O(N__5752),
            .I(Gl_r2_2));
    Odrv4 I__1229 (
            .O(N__5749),
            .I(Gl_r2_2));
    InMux I__1228 (
            .O(N__5734),
            .I(N__5728));
    InMux I__1227 (
            .O(N__5733),
            .I(N__5728));
    LocalMux I__1226 (
            .O(N__5728),
            .I(N__5725));
    Span4Mux_h I__1225 (
            .O(N__5725),
            .I(N__5712));
    InMux I__1224 (
            .O(N__5724),
            .I(N__5707));
    InMux I__1223 (
            .O(N__5723),
            .I(N__5707));
    InMux I__1222 (
            .O(N__5722),
            .I(N__5702));
    InMux I__1221 (
            .O(N__5721),
            .I(N__5702));
    InMux I__1220 (
            .O(N__5720),
            .I(N__5695));
    InMux I__1219 (
            .O(N__5719),
            .I(N__5695));
    InMux I__1218 (
            .O(N__5718),
            .I(N__5695));
    InMux I__1217 (
            .O(N__5717),
            .I(N__5688));
    InMux I__1216 (
            .O(N__5716),
            .I(N__5688));
    InMux I__1215 (
            .O(N__5715),
            .I(N__5688));
    Odrv4 I__1214 (
            .O(N__5712),
            .I(Gl_r1_3));
    LocalMux I__1213 (
            .O(N__5707),
            .I(Gl_r1_3));
    LocalMux I__1212 (
            .O(N__5702),
            .I(Gl_r1_3));
    LocalMux I__1211 (
            .O(N__5695),
            .I(Gl_r1_3));
    LocalMux I__1210 (
            .O(N__5688),
            .I(Gl_r1_3));
    InMux I__1209 (
            .O(N__5677),
            .I(N__5674));
    LocalMux I__1208 (
            .O(N__5674),
            .I(N__5671));
    Span4Mux_v I__1207 (
            .O(N__5671),
            .I(N__5668));
    Odrv4 I__1206 (
            .O(N__5668),
            .I(\Lab_UT.S_1_c3_d ));
    CascadeMux I__1205 (
            .O(N__5665),
            .I(\Lab_UT.S_1_c3_cZ0_cascade_ ));
    CascadeMux I__1204 (
            .O(N__5662),
            .I(N__5657));
    CascadeMux I__1203 (
            .O(N__5661),
            .I(N__5653));
    InMux I__1202 (
            .O(N__5660),
            .I(N__5646));
    InMux I__1201 (
            .O(N__5657),
            .I(N__5646));
    CascadeMux I__1200 (
            .O(N__5656),
            .I(N__5643));
    InMux I__1199 (
            .O(N__5653),
            .I(N__5634));
    InMux I__1198 (
            .O(N__5652),
            .I(N__5634));
    InMux I__1197 (
            .O(N__5651),
            .I(N__5634));
    LocalMux I__1196 (
            .O(N__5646),
            .I(N__5627));
    InMux I__1195 (
            .O(N__5643),
            .I(N__5620));
    InMux I__1194 (
            .O(N__5642),
            .I(N__5620));
    InMux I__1193 (
            .O(N__5641),
            .I(N__5620));
    LocalMux I__1192 (
            .O(N__5634),
            .I(N__5617));
    InMux I__1191 (
            .O(N__5633),
            .I(N__5612));
    InMux I__1190 (
            .O(N__5632),
            .I(N__5612));
    InMux I__1189 (
            .O(N__5631),
            .I(N__5607));
    InMux I__1188 (
            .O(N__5630),
            .I(N__5607));
    Span4Mux_h I__1187 (
            .O(N__5627),
            .I(N__5602));
    LocalMux I__1186 (
            .O(N__5620),
            .I(N__5602));
    Odrv4 I__1185 (
            .O(N__5617),
            .I(Gl_r2_3));
    LocalMux I__1184 (
            .O(N__5612),
            .I(Gl_r2_3));
    LocalMux I__1183 (
            .O(N__5607),
            .I(Gl_r2_3));
    Odrv4 I__1182 (
            .O(N__5602),
            .I(Gl_r2_3));
    InMux I__1181 (
            .O(N__5593),
            .I(N__5590));
    LocalMux I__1180 (
            .O(N__5590),
            .I(\Lab_UT.S_0_s_ac0_5_0Z0Z_0 ));
    InMux I__1179 (
            .O(N__5587),
            .I(N__5584));
    LocalMux I__1178 (
            .O(N__5584),
            .I(N__5581));
    Span4Mux_v I__1177 (
            .O(N__5581),
            .I(N__5578));
    Odrv4 I__1176 (
            .O(N__5578),
            .I(\Lab_UT.S_0_s_ac0_5_dZ0 ));
    CascadeMux I__1175 (
            .O(N__5575),
            .I(\Lab_UT.C_out41_cascade_ ));
    InMux I__1174 (
            .O(N__5572),
            .I(N__5568));
    InMux I__1173 (
            .O(N__5571),
            .I(N__5565));
    LocalMux I__1172 (
            .O(N__5568),
            .I(N__5562));
    LocalMux I__1171 (
            .O(N__5565),
            .I(N__5559));
    Span4Mux_s3_h I__1170 (
            .O(N__5562),
            .I(N__5552));
    Span4Mux_h I__1169 (
            .O(N__5559),
            .I(N__5552));
    InMux I__1168 (
            .O(N__5558),
            .I(N__5547));
    InMux I__1167 (
            .O(N__5557),
            .I(N__5547));
    Odrv4 I__1166 (
            .O(N__5552),
            .I(Gl_subtract));
    LocalMux I__1165 (
            .O(N__5547),
            .I(Gl_subtract));
    IoInMux I__1164 (
            .O(N__5542),
            .I(N__5539));
    LocalMux I__1163 (
            .O(N__5539),
            .I(N__5536));
    Span4Mux_s2_h I__1162 (
            .O(N__5536),
            .I(N__5533));
    Span4Mux_v I__1161 (
            .O(N__5533),
            .I(N__5530));
    Odrv4 I__1160 (
            .O(N__5530),
            .I(led_c_4));
    CascadeMux I__1159 (
            .O(N__5527),
            .I(\Glue_Lab2.de0.g0_5_1_cascade_ ));
    CascadeMux I__1158 (
            .O(N__5524),
            .I(\Glue_Lab2.g0_9_1_cascade_ ));
    InMux I__1157 (
            .O(N__5521),
            .I(N__5518));
    LocalMux I__1156 (
            .O(N__5518),
            .I(N__5515));
    Span4Mux_v I__1155 (
            .O(N__5515),
            .I(N__5512));
    Odrv4 I__1154 (
            .O(N__5512),
            .I(\Glue_Lab2.g0_7_1 ));
    InMux I__1153 (
            .O(N__5509),
            .I(N__5506));
    LocalMux I__1152 (
            .O(N__5506),
            .I(N__5503));
    Odrv12 I__1151 (
            .O(N__5503),
            .I(\Glue_Lab2.reset_counte_0_2 ));
    InMux I__1150 (
            .O(N__5500),
            .I(N__5496));
    InMux I__1149 (
            .O(N__5499),
            .I(N__5490));
    LocalMux I__1148 (
            .O(N__5496),
            .I(N__5484));
    InMux I__1147 (
            .O(N__5495),
            .I(N__5477));
    InMux I__1146 (
            .O(N__5494),
            .I(N__5477));
    InMux I__1145 (
            .O(N__5493),
            .I(N__5477));
    LocalMux I__1144 (
            .O(N__5490),
            .I(N__5474));
    InMux I__1143 (
            .O(N__5489),
            .I(N__5467));
    InMux I__1142 (
            .O(N__5488),
            .I(N__5467));
    InMux I__1141 (
            .O(N__5487),
            .I(N__5467));
    Span4Mux_v I__1140 (
            .O(N__5484),
            .I(N__5462));
    LocalMux I__1139 (
            .O(N__5477),
            .I(N__5462));
    Odrv4 I__1138 (
            .O(N__5474),
            .I(bu_rx_data_4));
    LocalMux I__1137 (
            .O(N__5467),
            .I(bu_rx_data_4));
    Odrv4 I__1136 (
            .O(N__5462),
            .I(bu_rx_data_4));
    InMux I__1135 (
            .O(N__5455),
            .I(N__5448));
    InMux I__1134 (
            .O(N__5454),
            .I(N__5448));
    InMux I__1133 (
            .O(N__5453),
            .I(N__5444));
    LocalMux I__1132 (
            .O(N__5448),
            .I(N__5440));
    InMux I__1131 (
            .O(N__5447),
            .I(N__5432));
    LocalMux I__1130 (
            .O(N__5444),
            .I(N__5429));
    InMux I__1129 (
            .O(N__5443),
            .I(N__5426));
    Span4Mux_s3_h I__1128 (
            .O(N__5440),
            .I(N__5423));
    InMux I__1127 (
            .O(N__5439),
            .I(N__5420));
    InMux I__1126 (
            .O(N__5438),
            .I(N__5417));
    InMux I__1125 (
            .O(N__5437),
            .I(N__5414));
    InMux I__1124 (
            .O(N__5436),
            .I(N__5409));
    InMux I__1123 (
            .O(N__5435),
            .I(N__5409));
    LocalMux I__1122 (
            .O(N__5432),
            .I(buart__rx_bitcount_0));
    Odrv4 I__1121 (
            .O(N__5429),
            .I(buart__rx_bitcount_0));
    LocalMux I__1120 (
            .O(N__5426),
            .I(buart__rx_bitcount_0));
    Odrv4 I__1119 (
            .O(N__5423),
            .I(buart__rx_bitcount_0));
    LocalMux I__1118 (
            .O(N__5420),
            .I(buart__rx_bitcount_0));
    LocalMux I__1117 (
            .O(N__5417),
            .I(buart__rx_bitcount_0));
    LocalMux I__1116 (
            .O(N__5414),
            .I(buart__rx_bitcount_0));
    LocalMux I__1115 (
            .O(N__5409),
            .I(buart__rx_bitcount_0));
    CascadeMux I__1114 (
            .O(N__5392),
            .I(\Glue_Lab2.de0.g0Z0Z_5_cascade_ ));
    InMux I__1113 (
            .O(N__5389),
            .I(N__5377));
    InMux I__1112 (
            .O(N__5388),
            .I(N__5377));
    InMux I__1111 (
            .O(N__5387),
            .I(N__5374));
    InMux I__1110 (
            .O(N__5386),
            .I(N__5371));
    InMux I__1109 (
            .O(N__5385),
            .I(N__5366));
    InMux I__1108 (
            .O(N__5384),
            .I(N__5366));
    InMux I__1107 (
            .O(N__5383),
            .I(N__5363));
    InMux I__1106 (
            .O(N__5382),
            .I(N__5360));
    LocalMux I__1105 (
            .O(N__5377),
            .I(N__5357));
    LocalMux I__1104 (
            .O(N__5374),
            .I(N__5352));
    LocalMux I__1103 (
            .O(N__5371),
            .I(N__5349));
    LocalMux I__1102 (
            .O(N__5366),
            .I(N__5346));
    LocalMux I__1101 (
            .O(N__5363),
            .I(N__5341));
    LocalMux I__1100 (
            .O(N__5360),
            .I(N__5336));
    Span4Mux_v I__1099 (
            .O(N__5357),
            .I(N__5336));
    InMux I__1098 (
            .O(N__5356),
            .I(N__5331));
    InMux I__1097 (
            .O(N__5355),
            .I(N__5331));
    Span4Mux_h I__1096 (
            .O(N__5352),
            .I(N__5328));
    Span4Mux_h I__1095 (
            .O(N__5349),
            .I(N__5323));
    Span4Mux_s2_h I__1094 (
            .O(N__5346),
            .I(N__5323));
    InMux I__1093 (
            .O(N__5345),
            .I(N__5318));
    InMux I__1092 (
            .O(N__5344),
            .I(N__5318));
    Odrv4 I__1091 (
            .O(N__5341),
            .I(bu_rx_data_0));
    Odrv4 I__1090 (
            .O(N__5336),
            .I(bu_rx_data_0));
    LocalMux I__1089 (
            .O(N__5331),
            .I(bu_rx_data_0));
    Odrv4 I__1088 (
            .O(N__5328),
            .I(bu_rx_data_0));
    Odrv4 I__1087 (
            .O(N__5323),
            .I(bu_rx_data_0));
    LocalMux I__1086 (
            .O(N__5318),
            .I(bu_rx_data_0));
    InMux I__1085 (
            .O(N__5305),
            .I(N__5300));
    InMux I__1084 (
            .O(N__5304),
            .I(N__5295));
    InMux I__1083 (
            .O(N__5303),
            .I(N__5295));
    LocalMux I__1082 (
            .O(N__5300),
            .I(N__5289));
    LocalMux I__1081 (
            .O(N__5295),
            .I(N__5286));
    InMux I__1080 (
            .O(N__5294),
            .I(N__5283));
    InMux I__1079 (
            .O(N__5293),
            .I(N__5280));
    InMux I__1078 (
            .O(N__5292),
            .I(N__5277));
    Span4Mux_h I__1077 (
            .O(N__5289),
            .I(N__5274));
    Span4Mux_s2_h I__1076 (
            .O(N__5286),
            .I(N__5269));
    LocalMux I__1075 (
            .O(N__5283),
            .I(N__5269));
    LocalMux I__1074 (
            .O(N__5280),
            .I(\Glue_Lab2.reset_countZ0Z_4 ));
    LocalMux I__1073 (
            .O(N__5277),
            .I(\Glue_Lab2.reset_countZ0Z_4 ));
    Odrv4 I__1072 (
            .O(N__5274),
            .I(\Glue_Lab2.reset_countZ0Z_4 ));
    Odrv4 I__1071 (
            .O(N__5269),
            .I(\Glue_Lab2.reset_countZ0Z_4 ));
    CascadeMux I__1070 (
            .O(N__5260),
            .I(\Glue_Lab2.g0_9_cascade_ ));
    InMux I__1069 (
            .O(N__5257),
            .I(N__5254));
    LocalMux I__1068 (
            .O(N__5254),
            .I(N__5251));
    Odrv4 I__1067 (
            .O(N__5251),
            .I(\Glue_Lab2.g0_7 ));
    InMux I__1066 (
            .O(N__5248),
            .I(N__5245));
    LocalMux I__1065 (
            .O(N__5245),
            .I(N__5242));
    Span4Mux_h I__1064 (
            .O(N__5242),
            .I(N__5239));
    Odrv4 I__1063 (
            .O(N__5239),
            .I(\Glue_Lab2.reset_counte_0_0 ));
    InMux I__1062 (
            .O(N__5236),
            .I(N__5223));
    InMux I__1061 (
            .O(N__5235),
            .I(N__5220));
    InMux I__1060 (
            .O(N__5234),
            .I(N__5213));
    InMux I__1059 (
            .O(N__5233),
            .I(N__5213));
    InMux I__1058 (
            .O(N__5232),
            .I(N__5213));
    InMux I__1057 (
            .O(N__5231),
            .I(N__5210));
    InMux I__1056 (
            .O(N__5230),
            .I(N__5207));
    InMux I__1055 (
            .O(N__5229),
            .I(N__5204));
    InMux I__1054 (
            .O(N__5228),
            .I(N__5201));
    InMux I__1053 (
            .O(N__5227),
            .I(N__5198));
    InMux I__1052 (
            .O(N__5226),
            .I(N__5193));
    LocalMux I__1051 (
            .O(N__5223),
            .I(N__5184));
    LocalMux I__1050 (
            .O(N__5220),
            .I(N__5184));
    LocalMux I__1049 (
            .O(N__5213),
            .I(N__5184));
    LocalMux I__1048 (
            .O(N__5210),
            .I(N__5184));
    LocalMux I__1047 (
            .O(N__5207),
            .I(N__5181));
    LocalMux I__1046 (
            .O(N__5204),
            .I(N__5178));
    LocalMux I__1045 (
            .O(N__5201),
            .I(N__5170));
    LocalMux I__1044 (
            .O(N__5198),
            .I(N__5170));
    InMux I__1043 (
            .O(N__5197),
            .I(N__5167));
    InMux I__1042 (
            .O(N__5196),
            .I(N__5164));
    LocalMux I__1041 (
            .O(N__5193),
            .I(N__5157));
    Span4Mux_v I__1040 (
            .O(N__5184),
            .I(N__5157));
    Span4Mux_v I__1039 (
            .O(N__5181),
            .I(N__5157));
    Span4Mux_h I__1038 (
            .O(N__5178),
            .I(N__5154));
    InMux I__1037 (
            .O(N__5177),
            .I(N__5147));
    InMux I__1036 (
            .O(N__5176),
            .I(N__5147));
    InMux I__1035 (
            .O(N__5175),
            .I(N__5147));
    Span12Mux_s4_v I__1034 (
            .O(N__5170),
            .I(N__5140));
    LocalMux I__1033 (
            .O(N__5167),
            .I(N__5140));
    LocalMux I__1032 (
            .O(N__5164),
            .I(N__5140));
    Odrv4 I__1031 (
            .O(N__5157),
            .I(bu_rx_data_2));
    Odrv4 I__1030 (
            .O(N__5154),
            .I(bu_rx_data_2));
    LocalMux I__1029 (
            .O(N__5147),
            .I(bu_rx_data_2));
    Odrv12 I__1028 (
            .O(N__5140),
            .I(bu_rx_data_2));
    InMux I__1027 (
            .O(N__5131),
            .I(N__5126));
    InMux I__1026 (
            .O(N__5130),
            .I(N__5123));
    CascadeMux I__1025 (
            .O(N__5129),
            .I(N__5120));
    LocalMux I__1024 (
            .O(N__5126),
            .I(N__5115));
    LocalMux I__1023 (
            .O(N__5123),
            .I(N__5112));
    InMux I__1022 (
            .O(N__5120),
            .I(N__5105));
    InMux I__1021 (
            .O(N__5119),
            .I(N__5105));
    InMux I__1020 (
            .O(N__5118),
            .I(N__5105));
    Span4Mux_v I__1019 (
            .O(N__5115),
            .I(N__5092));
    Span4Mux_v I__1018 (
            .O(N__5112),
            .I(N__5092));
    LocalMux I__1017 (
            .O(N__5105),
            .I(N__5092));
    InMux I__1016 (
            .O(N__5104),
            .I(N__5089));
    InMux I__1015 (
            .O(N__5103),
            .I(N__5080));
    InMux I__1014 (
            .O(N__5102),
            .I(N__5080));
    InMux I__1013 (
            .O(N__5101),
            .I(N__5080));
    InMux I__1012 (
            .O(N__5100),
            .I(N__5080));
    InMux I__1011 (
            .O(N__5099),
            .I(N__5077));
    Odrv4 I__1010 (
            .O(N__5092),
            .I(bu_rx_data_6));
    LocalMux I__1009 (
            .O(N__5089),
            .I(bu_rx_data_6));
    LocalMux I__1008 (
            .O(N__5080),
            .I(bu_rx_data_6));
    LocalMux I__1007 (
            .O(N__5077),
            .I(bu_rx_data_6));
    InMux I__1006 (
            .O(N__5068),
            .I(N__5059));
    InMux I__1005 (
            .O(N__5067),
            .I(N__5059));
    InMux I__1004 (
            .O(N__5066),
            .I(N__5059));
    LocalMux I__1003 (
            .O(N__5059),
            .I(\buart.Z_tx.bitcountZ0Z_2 ));
    CascadeMux I__1002 (
            .O(N__5056),
            .I(\buart.Z_tx.un1_bitcount_c3_cascade_ ));
    InMux I__1001 (
            .O(N__5053),
            .I(N__5047));
    InMux I__1000 (
            .O(N__5052),
            .I(N__5047));
    LocalMux I__999 (
            .O(N__5047),
            .I(\buart.Z_tx.bitcountZ0Z_3 ));
    InMux I__998 (
            .O(N__5044),
            .I(N__5041));
    LocalMux I__997 (
            .O(N__5041),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i_sx ));
    InMux I__996 (
            .O(N__5038),
            .I(N__5034));
    CascadeMux I__995 (
            .O(N__5037),
            .I(N__5028));
    LocalMux I__994 (
            .O(N__5034),
            .I(N__5025));
    InMux I__993 (
            .O(N__5033),
            .I(N__5022));
    InMux I__992 (
            .O(N__5032),
            .I(N__5019));
    InMux I__991 (
            .O(N__5031),
            .I(N__5011));
    InMux I__990 (
            .O(N__5028),
            .I(N__5011));
    Span4Mux_s3_h I__989 (
            .O(N__5025),
            .I(N__5005));
    LocalMux I__988 (
            .O(N__5022),
            .I(N__5000));
    LocalMux I__987 (
            .O(N__5019),
            .I(N__5000));
    InMux I__986 (
            .O(N__5018),
            .I(N__4995));
    InMux I__985 (
            .O(N__5017),
            .I(N__4995));
    InMux I__984 (
            .O(N__5016),
            .I(N__4992));
    LocalMux I__983 (
            .O(N__5011),
            .I(N__4989));
    InMux I__982 (
            .O(N__5010),
            .I(N__4982));
    InMux I__981 (
            .O(N__5009),
            .I(N__4982));
    InMux I__980 (
            .O(N__5008),
            .I(N__4982));
    Odrv4 I__979 (
            .O(N__5005),
            .I(\Glue_Lab2.is_hexplus ));
    Odrv4 I__978 (
            .O(N__5000),
            .I(\Glue_Lab2.is_hexplus ));
    LocalMux I__977 (
            .O(N__4995),
            .I(\Glue_Lab2.is_hexplus ));
    LocalMux I__976 (
            .O(N__4992),
            .I(\Glue_Lab2.is_hexplus ));
    Odrv4 I__975 (
            .O(N__4989),
            .I(\Glue_Lab2.is_hexplus ));
    LocalMux I__974 (
            .O(N__4982),
            .I(\Glue_Lab2.is_hexplus ));
    CascadeMux I__973 (
            .O(N__4969),
            .I(\buart.Z_tx.un1_bitcount_c1_cascade_ ));
    CascadeMux I__972 (
            .O(N__4966),
            .I(N__4962));
    InMux I__971 (
            .O(N__4965),
            .I(N__4956));
    InMux I__970 (
            .O(N__4962),
            .I(N__4949));
    InMux I__969 (
            .O(N__4961),
            .I(N__4949));
    InMux I__968 (
            .O(N__4960),
            .I(N__4949));
    InMux I__967 (
            .O(N__4959),
            .I(N__4946));
    LocalMux I__966 (
            .O(N__4956),
            .I(\buart.Z_tx.bitcountZ0Z_1 ));
    LocalMux I__965 (
            .O(N__4949),
            .I(\buart.Z_tx.bitcountZ0Z_1 ));
    LocalMux I__964 (
            .O(N__4946),
            .I(\buart.Z_tx.bitcountZ0Z_1 ));
    InMux I__963 (
            .O(N__4939),
            .I(N__4934));
    InMux I__962 (
            .O(N__4938),
            .I(N__4929));
    InMux I__961 (
            .O(N__4937),
            .I(N__4929));
    LocalMux I__960 (
            .O(N__4934),
            .I(\buart.Z_tx.counter_RNIVE1P1_4 ));
    LocalMux I__959 (
            .O(N__4929),
            .I(\buart.Z_tx.counter_RNIVE1P1_4 ));
    InMux I__958 (
            .O(N__4924),
            .I(N__4914));
    InMux I__957 (
            .O(N__4923),
            .I(N__4914));
    InMux I__956 (
            .O(N__4922),
            .I(N__4905));
    InMux I__955 (
            .O(N__4921),
            .I(N__4905));
    InMux I__954 (
            .O(N__4920),
            .I(N__4905));
    InMux I__953 (
            .O(N__4919),
            .I(N__4905));
    LocalMux I__952 (
            .O(N__4914),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    LocalMux I__951 (
            .O(N__4905),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    InMux I__950 (
            .O(N__4900),
            .I(N__4897));
    LocalMux I__949 (
            .O(N__4897),
            .I(N__4894));
    Span4Mux_h I__948 (
            .O(N__4894),
            .I(N__4891));
    Odrv4 I__947 (
            .O(N__4891),
            .I(\Glue_Lab2.de0.de_escZ0Z_4 ));
    InMux I__946 (
            .O(N__4888),
            .I(N__4876));
    InMux I__945 (
            .O(N__4887),
            .I(N__4876));
    InMux I__944 (
            .O(N__4886),
            .I(N__4876));
    InMux I__943 (
            .O(N__4885),
            .I(N__4876));
    LocalMux I__942 (
            .O(N__4876),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ));
    CascadeMux I__941 (
            .O(N__4873),
            .I(N__4867));
    InMux I__940 (
            .O(N__4872),
            .I(N__4858));
    InMux I__939 (
            .O(N__4871),
            .I(N__4858));
    InMux I__938 (
            .O(N__4870),
            .I(N__4858));
    InMux I__937 (
            .O(N__4867),
            .I(N__4858));
    LocalMux I__936 (
            .O(N__4858),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_5 ));
    InMux I__935 (
            .O(N__4855),
            .I(N__4846));
    InMux I__934 (
            .O(N__4854),
            .I(N__4846));
    InMux I__933 (
            .O(N__4853),
            .I(N__4846));
    LocalMux I__932 (
            .O(N__4846),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ));
    CascadeMux I__931 (
            .O(N__4843),
            .I(N__4840));
    InMux I__930 (
            .O(N__4840),
            .I(N__4832));
    InMux I__929 (
            .O(N__4839),
            .I(N__4832));
    InMux I__928 (
            .O(N__4838),
            .I(N__4827));
    InMux I__927 (
            .O(N__4837),
            .I(N__4827));
    LocalMux I__926 (
            .O(N__4832),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    LocalMux I__925 (
            .O(N__4827),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    CascadeMux I__924 (
            .O(N__4822),
            .I(\buart.Z_tx.Z_baudgen.ser_clk_sx_cascade_ ));
    InMux I__923 (
            .O(N__4819),
            .I(N__4808));
    InMux I__922 (
            .O(N__4818),
            .I(N__4808));
    InMux I__921 (
            .O(N__4817),
            .I(N__4808));
    InMux I__920 (
            .O(N__4816),
            .I(N__4803));
    InMux I__919 (
            .O(N__4815),
            .I(N__4803));
    LocalMux I__918 (
            .O(N__4808),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__917 (
            .O(N__4803),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    InMux I__916 (
            .O(N__4798),
            .I(N__4795));
    LocalMux I__915 (
            .O(N__4795),
            .I(\buart.Z_tx.Z_baudgen.counter_RNIES38_0Z0Z_4 ));
    InMux I__914 (
            .O(N__4792),
            .I(N__4789));
    LocalMux I__913 (
            .O(N__4789),
            .I(\buart.Z_tx.Z_baudgen.un1_bitcount_c2_1 ));
    CascadeMux I__912 (
            .O(N__4786),
            .I(\buart.Z_tx.bitcount_RNIBADLZ0Z_1_cascade_ ));
    CascadeMux I__911 (
            .O(N__4783),
            .I(\buart.Z_tx.counter_RNIVE1P1_4_cascade_ ));
    InMux I__910 (
            .O(N__4780),
            .I(N__4777));
    LocalMux I__909 (
            .O(N__4777),
            .I(\buart.Z_tx.un1_bitcount_c2 ));
    InMux I__908 (
            .O(N__4774),
            .I(N__4771));
    LocalMux I__907 (
            .O(N__4771),
            .I(\buart.Z_tx.uart_busy_0_0 ));
    CascadeMux I__906 (
            .O(N__4768),
            .I(\buart.Z_tx.uart_busy_0_0_cascade_ ));
    CascadeMux I__905 (
            .O(N__4765),
            .I(led_c_1_cascade_));
    InMux I__904 (
            .O(N__4762),
            .I(N__4759));
    LocalMux I__903 (
            .O(N__4759),
            .I(N__4756));
    Span12Mux_s8_h I__902 (
            .O(N__4756),
            .I(N__4753));
    Odrv12 I__901 (
            .O(N__4753),
            .I(Gl_tx_data_1));
    InMux I__900 (
            .O(N__4750),
            .I(N__4747));
    LocalMux I__899 (
            .O(N__4747),
            .I(N__4743));
    InMux I__898 (
            .O(N__4746),
            .I(N__4740));
    Odrv4 I__897 (
            .O(N__4743),
            .I(Gl_r2_fast_2));
    LocalMux I__896 (
            .O(N__4740),
            .I(Gl_r2_fast_2));
    InMux I__895 (
            .O(N__4735),
            .I(N__4731));
    InMux I__894 (
            .O(N__4734),
            .I(N__4728));
    LocalMux I__893 (
            .O(N__4731),
            .I(Gl_r1_fast_2));
    LocalMux I__892 (
            .O(N__4728),
            .I(Gl_r1_fast_2));
    InMux I__891 (
            .O(N__4723),
            .I(N__4720));
    LocalMux I__890 (
            .O(N__4720),
            .I(\Lab_UT.S_m_bm_1Z0Z_2 ));
    InMux I__889 (
            .O(N__4717),
            .I(N__4714));
    LocalMux I__888 (
            .O(N__4714),
            .I(\Lab_UT.S_m_bmZ0Z_2 ));
    CascadeMux I__887 (
            .O(N__4711),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_c5_cascade_ ));
    CascadeMux I__886 (
            .O(N__4708),
            .I(N__4705));
    InMux I__885 (
            .O(N__4705),
            .I(N__4702));
    LocalMux I__884 (
            .O(N__4702),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_c5 ));
    InMux I__883 (
            .O(N__4699),
            .I(N__4690));
    InMux I__882 (
            .O(N__4698),
            .I(N__4690));
    InMux I__881 (
            .O(N__4697),
            .I(N__4686));
    InMux I__880 (
            .O(N__4696),
            .I(N__4681));
    InMux I__879 (
            .O(N__4695),
            .I(N__4681));
    LocalMux I__878 (
            .O(N__4690),
            .I(N__4678));
    InMux I__877 (
            .O(N__4689),
            .I(N__4675));
    LocalMux I__876 (
            .O(N__4686),
            .I(Glue_Lab2_gl_fsm_state_1));
    LocalMux I__875 (
            .O(N__4681),
            .I(Glue_Lab2_gl_fsm_state_1));
    Odrv4 I__874 (
            .O(N__4678),
            .I(Glue_Lab2_gl_fsm_state_1));
    LocalMux I__873 (
            .O(N__4675),
            .I(Glue_Lab2_gl_fsm_state_1));
    InMux I__872 (
            .O(N__4666),
            .I(N__4663));
    LocalMux I__871 (
            .O(N__4663),
            .I(N__4660));
    Odrv4 I__870 (
            .O(N__4660),
            .I(\Glue_Lab2.gl_fsm.enOp_0_a2_2 ));
    CascadeMux I__869 (
            .O(N__4657),
            .I(\Glue_Lab2.Gl_subtract_1_cascade_ ));
    InMux I__868 (
            .O(N__4654),
            .I(N__4651));
    LocalMux I__867 (
            .O(N__4651),
            .I(N__4648));
    Odrv12 I__866 (
            .O(N__4648),
            .I(\Lab_UT.S_0_s_axbZ0Z3 ));
    CascadeMux I__865 (
            .O(N__4645),
            .I(N__4642));
    InMux I__864 (
            .O(N__4642),
            .I(N__4636));
    InMux I__863 (
            .O(N__4641),
            .I(N__4636));
    LocalMux I__862 (
            .O(N__4636),
            .I(N__4632));
    InMux I__861 (
            .O(N__4635),
            .I(N__4629));
    Odrv4 I__860 (
            .O(N__4632),
            .I(\Lab_UT.S_0_s_cZ0Z2 ));
    LocalMux I__859 (
            .O(N__4629),
            .I(\Lab_UT.S_0_s_cZ0Z2 ));
    CascadeMux I__858 (
            .O(N__4624),
            .I(\Lab_UT.S_m_amZ0Z_2_cascade_ ));
    IoInMux I__857 (
            .O(N__4621),
            .I(N__4618));
    LocalMux I__856 (
            .O(N__4618),
            .I(N__4615));
    Span4Mux_s3_h I__855 (
            .O(N__4615),
            .I(N__4611));
    InMux I__854 (
            .O(N__4614),
            .I(N__4608));
    Odrv4 I__853 (
            .O(N__4611),
            .I(led_c_2));
    LocalMux I__852 (
            .O(N__4608),
            .I(led_c_2));
    InMux I__851 (
            .O(N__4603),
            .I(N__4598));
    CascadeMux I__850 (
            .O(N__4602),
            .I(N__4591));
    InMux I__849 (
            .O(N__4601),
            .I(N__4587));
    LocalMux I__848 (
            .O(N__4598),
            .I(N__4584));
    InMux I__847 (
            .O(N__4597),
            .I(N__4581));
    InMux I__846 (
            .O(N__4596),
            .I(N__4578));
    InMux I__845 (
            .O(N__4595),
            .I(N__4569));
    InMux I__844 (
            .O(N__4594),
            .I(N__4569));
    InMux I__843 (
            .O(N__4591),
            .I(N__4569));
    InMux I__842 (
            .O(N__4590),
            .I(N__4569));
    LocalMux I__841 (
            .O(N__4587),
            .I(Gl_r1_0));
    Odrv4 I__840 (
            .O(N__4584),
            .I(Gl_r1_0));
    LocalMux I__839 (
            .O(N__4581),
            .I(Gl_r1_0));
    LocalMux I__838 (
            .O(N__4578),
            .I(Gl_r1_0));
    LocalMux I__837 (
            .O(N__4569),
            .I(Gl_r1_0));
    CascadeMux I__836 (
            .O(N__4558),
            .I(N__4553));
    CascadeMux I__835 (
            .O(N__4557),
            .I(N__4543));
    InMux I__834 (
            .O(N__4556),
            .I(N__4532));
    InMux I__833 (
            .O(N__4553),
            .I(N__4532));
    InMux I__832 (
            .O(N__4552),
            .I(N__4532));
    InMux I__831 (
            .O(N__4551),
            .I(N__4532));
    InMux I__830 (
            .O(N__4550),
            .I(N__4532));
    InMux I__829 (
            .O(N__4549),
            .I(N__4529));
    InMux I__828 (
            .O(N__4548),
            .I(N__4523));
    InMux I__827 (
            .O(N__4547),
            .I(N__4520));
    InMux I__826 (
            .O(N__4546),
            .I(N__4515));
    InMux I__825 (
            .O(N__4543),
            .I(N__4515));
    LocalMux I__824 (
            .O(N__4532),
            .I(N__4510));
    LocalMux I__823 (
            .O(N__4529),
            .I(N__4510));
    InMux I__822 (
            .O(N__4528),
            .I(N__4505));
    InMux I__821 (
            .O(N__4527),
            .I(N__4505));
    InMux I__820 (
            .O(N__4526),
            .I(N__4502));
    LocalMux I__819 (
            .O(N__4523),
            .I(Gl_r2_1));
    LocalMux I__818 (
            .O(N__4520),
            .I(Gl_r2_1));
    LocalMux I__817 (
            .O(N__4515),
            .I(Gl_r2_1));
    Odrv4 I__816 (
            .O(N__4510),
            .I(Gl_r2_1));
    LocalMux I__815 (
            .O(N__4505),
            .I(Gl_r2_1));
    LocalMux I__814 (
            .O(N__4502),
            .I(Gl_r2_1));
    CascadeMux I__813 (
            .O(N__4489),
            .I(N__4482));
    CascadeMux I__812 (
            .O(N__4488),
            .I(N__4479));
    CascadeMux I__811 (
            .O(N__4487),
            .I(N__4475));
    CascadeMux I__810 (
            .O(N__4486),
            .I(N__4471));
    InMux I__809 (
            .O(N__4485),
            .I(N__4468));
    InMux I__808 (
            .O(N__4482),
            .I(N__4465));
    InMux I__807 (
            .O(N__4479),
            .I(N__4462));
    InMux I__806 (
            .O(N__4478),
            .I(N__4453));
    InMux I__805 (
            .O(N__4475),
            .I(N__4453));
    InMux I__804 (
            .O(N__4474),
            .I(N__4453));
    InMux I__803 (
            .O(N__4471),
            .I(N__4453));
    LocalMux I__802 (
            .O(N__4468),
            .I(N__4450));
    LocalMux I__801 (
            .O(N__4465),
            .I(N__4444));
    LocalMux I__800 (
            .O(N__4462),
            .I(N__4444));
    LocalMux I__799 (
            .O(N__4453),
            .I(N__4441));
    Span4Mux_v I__798 (
            .O(N__4450),
            .I(N__4438));
    InMux I__797 (
            .O(N__4449),
            .I(N__4435));
    Span4Mux_h I__796 (
            .O(N__4444),
            .I(N__4432));
    Span4Mux_h I__795 (
            .O(N__4441),
            .I(N__4429));
    Odrv4 I__794 (
            .O(N__4438),
            .I(Gl_r2_0));
    LocalMux I__793 (
            .O(N__4435),
            .I(Gl_r2_0));
    Odrv4 I__792 (
            .O(N__4432),
            .I(Gl_r2_0));
    Odrv4 I__791 (
            .O(N__4429),
            .I(Gl_r2_0));
    InMux I__790 (
            .O(N__4420),
            .I(N__4417));
    LocalMux I__789 (
            .O(N__4417),
            .I(N__4411));
    InMux I__788 (
            .O(N__4416),
            .I(N__4406));
    InMux I__787 (
            .O(N__4415),
            .I(N__4406));
    CascadeMux I__786 (
            .O(N__4414),
            .I(N__4403));
    Span4Mux_s2_v I__785 (
            .O(N__4411),
            .I(N__4391));
    LocalMux I__784 (
            .O(N__4406),
            .I(N__4388));
    InMux I__783 (
            .O(N__4403),
            .I(N__4385));
    InMux I__782 (
            .O(N__4402),
            .I(N__4374));
    InMux I__781 (
            .O(N__4401),
            .I(N__4374));
    InMux I__780 (
            .O(N__4400),
            .I(N__4374));
    InMux I__779 (
            .O(N__4399),
            .I(N__4374));
    InMux I__778 (
            .O(N__4398),
            .I(N__4374));
    InMux I__777 (
            .O(N__4397),
            .I(N__4367));
    InMux I__776 (
            .O(N__4396),
            .I(N__4367));
    InMux I__775 (
            .O(N__4395),
            .I(N__4367));
    InMux I__774 (
            .O(N__4394),
            .I(N__4364));
    Odrv4 I__773 (
            .O(N__4391),
            .I(Gl_r1_1));
    Odrv4 I__772 (
            .O(N__4388),
            .I(Gl_r1_1));
    LocalMux I__771 (
            .O(N__4385),
            .I(Gl_r1_1));
    LocalMux I__770 (
            .O(N__4374),
            .I(Gl_r1_1));
    LocalMux I__769 (
            .O(N__4367),
            .I(Gl_r1_1));
    LocalMux I__768 (
            .O(N__4364),
            .I(Gl_r1_1));
    InMux I__767 (
            .O(N__4351),
            .I(N__4348));
    LocalMux I__766 (
            .O(N__4348),
            .I(\Lab_UT.S_m_amZ0Z_1 ));
    CascadeMux I__765 (
            .O(N__4345),
            .I(\Lab_UT.S_m_bmZ0Z_1_cascade_ ));
    IoInMux I__764 (
            .O(N__4342),
            .I(N__4339));
    LocalMux I__763 (
            .O(N__4339),
            .I(N__4336));
    Span4Mux_s3_h I__762 (
            .O(N__4336),
            .I(N__4333));
    Odrv4 I__761 (
            .O(N__4333),
            .I(led_c_1));
    InMux I__760 (
            .O(N__4330),
            .I(N__4327));
    LocalMux I__759 (
            .O(N__4327),
            .I(\Glue_Lab2.gl_fsm.enOp_0_a2_1 ));
    CascadeMux I__758 (
            .O(N__4324),
            .I(N__4321));
    InMux I__757 (
            .O(N__4321),
            .I(N__4318));
    LocalMux I__756 (
            .O(N__4318),
            .I(\Glue_Lab2.gl_fsm.enOp_0_a2Z0Z_4 ));
    InMux I__755 (
            .O(N__4315),
            .I(N__4309));
    InMux I__754 (
            .O(N__4314),
            .I(N__4304));
    InMux I__753 (
            .O(N__4313),
            .I(N__4304));
    InMux I__752 (
            .O(N__4312),
            .I(N__4301));
    LocalMux I__751 (
            .O(N__4309),
            .I(bu_rx_data_rdy));
    LocalMux I__750 (
            .O(N__4304),
            .I(bu_rx_data_rdy));
    LocalMux I__749 (
            .O(N__4301),
            .I(bu_rx_data_rdy));
    CascadeMux I__748 (
            .O(N__4294),
            .I(\Glue_Lab2.Gl_r1_2_1_cascade_ ));
    CascadeMux I__747 (
            .O(N__4291),
            .I(\Glue_Lab2.Gl_r1_2_2_cascade_ ));
    CascadeMux I__746 (
            .O(N__4288),
            .I(N__4285));
    InMux I__745 (
            .O(N__4285),
            .I(N__4282));
    LocalMux I__744 (
            .O(N__4282),
            .I(N__4279));
    Odrv4 I__743 (
            .O(N__4279),
            .I(\Lab_UT.g0Z0Z_1 ));
    CascadeMux I__742 (
            .O(N__4276),
            .I(N__4270));
    InMux I__741 (
            .O(N__4275),
            .I(N__4257));
    InMux I__740 (
            .O(N__4274),
            .I(N__4257));
    InMux I__739 (
            .O(N__4273),
            .I(N__4257));
    InMux I__738 (
            .O(N__4270),
            .I(N__4257));
    InMux I__737 (
            .O(N__4269),
            .I(N__4257));
    InMux I__736 (
            .O(N__4268),
            .I(N__4254));
    LocalMux I__735 (
            .O(N__4257),
            .I(\Glue_Lab2.enOp ));
    LocalMux I__734 (
            .O(N__4254),
            .I(\Glue_Lab2.enOp ));
    InMux I__733 (
            .O(N__4249),
            .I(N__4246));
    LocalMux I__732 (
            .O(N__4246),
            .I(N__4243));
    Span4Mux_h I__731 (
            .O(N__4243),
            .I(N__4240));
    Odrv4 I__730 (
            .O(N__4240),
            .I(Gl_tx_data_2));
    InMux I__729 (
            .O(N__4237),
            .I(N__4234));
    LocalMux I__728 (
            .O(N__4234),
            .I(\Glue_Lab2.de0.un1_charDataZ0 ));
    InMux I__727 (
            .O(N__4231),
            .I(N__4227));
    InMux I__726 (
            .O(N__4230),
            .I(N__4224));
    LocalMux I__725 (
            .O(N__4227),
            .I(buart__rx_shifter_fast_5));
    LocalMux I__724 (
            .O(N__4224),
            .I(buart__rx_shifter_fast_5));
    InMux I__723 (
            .O(N__4219),
            .I(N__4215));
    InMux I__722 (
            .O(N__4218),
            .I(N__4212));
    LocalMux I__721 (
            .O(N__4215),
            .I(N__4209));
    LocalMux I__720 (
            .O(N__4212),
            .I(N__4206));
    Span4Mux_v I__719 (
            .O(N__4209),
            .I(N__4201));
    Span4Mux_s3_h I__718 (
            .O(N__4206),
            .I(N__4201));
    Odrv4 I__717 (
            .O(N__4201),
            .I(\buart.Z_rx.hhZ0Z_1 ));
    InMux I__716 (
            .O(N__4198),
            .I(N__4195));
    LocalMux I__715 (
            .O(N__4195),
            .I(N__4192));
    Odrv4 I__714 (
            .O(N__4192),
            .I(\Glue_Lab2.g0_8_0 ));
    InMux I__713 (
            .O(N__4189),
            .I(N__4186));
    LocalMux I__712 (
            .O(N__4186),
            .I(\Glue_Lab2.de0.de_escZ0Z_3 ));
    CascadeMux I__711 (
            .O(N__4183),
            .I(N__4174));
    CascadeMux I__710 (
            .O(N__4182),
            .I(N__4171));
    CascadeMux I__709 (
            .O(N__4181),
            .I(N__4168));
    CascadeMux I__708 (
            .O(N__4180),
            .I(N__4165));
    CascadeMux I__707 (
            .O(N__4179),
            .I(N__4161));
    InMux I__706 (
            .O(N__4178),
            .I(N__4157));
    InMux I__705 (
            .O(N__4177),
            .I(N__4154));
    InMux I__704 (
            .O(N__4174),
            .I(N__4151));
    InMux I__703 (
            .O(N__4171),
            .I(N__4146));
    InMux I__702 (
            .O(N__4168),
            .I(N__4146));
    InMux I__701 (
            .O(N__4165),
            .I(N__4143));
    InMux I__700 (
            .O(N__4164),
            .I(N__4136));
    InMux I__699 (
            .O(N__4161),
            .I(N__4136));
    InMux I__698 (
            .O(N__4160),
            .I(N__4136));
    LocalMux I__697 (
            .O(N__4157),
            .I(buart__rx_bitcount_4));
    LocalMux I__696 (
            .O(N__4154),
            .I(buart__rx_bitcount_4));
    LocalMux I__695 (
            .O(N__4151),
            .I(buart__rx_bitcount_4));
    LocalMux I__694 (
            .O(N__4146),
            .I(buart__rx_bitcount_4));
    LocalMux I__693 (
            .O(N__4143),
            .I(buart__rx_bitcount_4));
    LocalMux I__692 (
            .O(N__4136),
            .I(buart__rx_bitcount_4));
    InMux I__691 (
            .O(N__4123),
            .I(N__4111));
    InMux I__690 (
            .O(N__4122),
            .I(N__4108));
    InMux I__689 (
            .O(N__4121),
            .I(N__4103));
    InMux I__688 (
            .O(N__4120),
            .I(N__4103));
    InMux I__687 (
            .O(N__4119),
            .I(N__4096));
    InMux I__686 (
            .O(N__4118),
            .I(N__4096));
    InMux I__685 (
            .O(N__4117),
            .I(N__4096));
    InMux I__684 (
            .O(N__4116),
            .I(N__4089));
    InMux I__683 (
            .O(N__4115),
            .I(N__4089));
    InMux I__682 (
            .O(N__4114),
            .I(N__4089));
    LocalMux I__681 (
            .O(N__4111),
            .I(buart__rx_bitcount_3));
    LocalMux I__680 (
            .O(N__4108),
            .I(buart__rx_bitcount_3));
    LocalMux I__679 (
            .O(N__4103),
            .I(buart__rx_bitcount_3));
    LocalMux I__678 (
            .O(N__4096),
            .I(buart__rx_bitcount_3));
    LocalMux I__677 (
            .O(N__4089),
            .I(buart__rx_bitcount_3));
    CascadeMux I__676 (
            .O(N__4078),
            .I(\buart.Z_rx.bitcount_RNIMK771Z0Z_4_cascade_ ));
    InMux I__675 (
            .O(N__4075),
            .I(N__4069));
    InMux I__674 (
            .O(N__4074),
            .I(N__4069));
    LocalMux I__673 (
            .O(N__4069),
            .I(\buart.Z_rx.idle ));
    CascadeMux I__672 (
            .O(N__4066),
            .I(\buart.Z_rx.idle_cascade_ ));
    InMux I__671 (
            .O(N__4063),
            .I(N__4060));
    LocalMux I__670 (
            .O(N__4060),
            .I(N__4056));
    InMux I__669 (
            .O(N__4059),
            .I(N__4053));
    Span4Mux_h I__668 (
            .O(N__4056),
            .I(N__4050));
    LocalMux I__667 (
            .O(N__4053),
            .I(\buart.Z_rx.hhZ0Z_0 ));
    Odrv4 I__666 (
            .O(N__4050),
            .I(\buart.Z_rx.hhZ0Z_0 ));
    CascadeMux I__665 (
            .O(N__4045),
            .I(\buart.Z_rx.startbit_cascade_ ));
    InMux I__664 (
            .O(N__4042),
            .I(N__4039));
    LocalMux I__663 (
            .O(N__4039),
            .I(\buart.Z_rx.bitcount_lm_1 ));
    InMux I__662 (
            .O(N__4036),
            .I(N__4022));
    InMux I__661 (
            .O(N__4035),
            .I(N__4022));
    InMux I__660 (
            .O(N__4034),
            .I(N__4015));
    InMux I__659 (
            .O(N__4033),
            .I(N__4015));
    InMux I__658 (
            .O(N__4032),
            .I(N__4015));
    InMux I__657 (
            .O(N__4031),
            .I(N__4010));
    InMux I__656 (
            .O(N__4030),
            .I(N__4010));
    InMux I__655 (
            .O(N__4029),
            .I(N__4003));
    InMux I__654 (
            .O(N__4028),
            .I(N__4003));
    InMux I__653 (
            .O(N__4027),
            .I(N__4003));
    LocalMux I__652 (
            .O(N__4022),
            .I(buart__rx_bitcount_1));
    LocalMux I__651 (
            .O(N__4015),
            .I(buart__rx_bitcount_1));
    LocalMux I__650 (
            .O(N__4010),
            .I(buart__rx_bitcount_1));
    LocalMux I__649 (
            .O(N__4003),
            .I(buart__rx_bitcount_1));
    InMux I__648 (
            .O(N__3994),
            .I(N__3991));
    LocalMux I__647 (
            .O(N__3991),
            .I(\buart.Z_rx.bitcount_cry_1_THRU_CO ));
    InMux I__646 (
            .O(N__3988),
            .I(N__3980));
    InMux I__645 (
            .O(N__3987),
            .I(N__3980));
    InMux I__644 (
            .O(N__3986),
            .I(N__3975));
    InMux I__643 (
            .O(N__3985),
            .I(N__3975));
    LocalMux I__642 (
            .O(N__3980),
            .I(\buart.Z_rx.N_29_0_i ));
    LocalMux I__641 (
            .O(N__3975),
            .I(\buart.Z_rx.N_29_0_i ));
    CascadeMux I__640 (
            .O(N__3970),
            .I(N__3964));
    InMux I__639 (
            .O(N__3969),
            .I(N__3957));
    InMux I__638 (
            .O(N__3968),
            .I(N__3957));
    InMux I__637 (
            .O(N__3967),
            .I(N__3957));
    InMux I__636 (
            .O(N__3964),
            .I(N__3954));
    LocalMux I__635 (
            .O(N__3957),
            .I(\buart.Z_rx.bitcountlde_0 ));
    LocalMux I__634 (
            .O(N__3954),
            .I(\buart.Z_rx.bitcountlde_0 ));
    CascadeMux I__633 (
            .O(N__3949),
            .I(\buart.Z_rx.bitcount_lm_2_cascade_ ));
    InMux I__632 (
            .O(N__3946),
            .I(N__3937));
    InMux I__631 (
            .O(N__3945),
            .I(N__3934));
    InMux I__630 (
            .O(N__3944),
            .I(N__3929));
    InMux I__629 (
            .O(N__3943),
            .I(N__3929));
    InMux I__628 (
            .O(N__3942),
            .I(N__3924));
    CascadeMux I__627 (
            .O(N__3941),
            .I(N__3919));
    CascadeMux I__626 (
            .O(N__3940),
            .I(N__3916));
    LocalMux I__625 (
            .O(N__3937),
            .I(N__3909));
    LocalMux I__624 (
            .O(N__3934),
            .I(N__3909));
    LocalMux I__623 (
            .O(N__3929),
            .I(N__3909));
    CascadeMux I__622 (
            .O(N__3928),
            .I(N__3902));
    CascadeMux I__621 (
            .O(N__3927),
            .I(N__3899));
    LocalMux I__620 (
            .O(N__3924),
            .I(N__3896));
    InMux I__619 (
            .O(N__3923),
            .I(N__3887));
    InMux I__618 (
            .O(N__3922),
            .I(N__3887));
    InMux I__617 (
            .O(N__3919),
            .I(N__3887));
    InMux I__616 (
            .O(N__3916),
            .I(N__3887));
    Span4Mux_v I__615 (
            .O(N__3909),
            .I(N__3884));
    InMux I__614 (
            .O(N__3908),
            .I(N__3875));
    InMux I__613 (
            .O(N__3907),
            .I(N__3875));
    InMux I__612 (
            .O(N__3906),
            .I(N__3875));
    InMux I__611 (
            .O(N__3905),
            .I(N__3875));
    InMux I__610 (
            .O(N__3902),
            .I(N__3872));
    InMux I__609 (
            .O(N__3899),
            .I(N__3869));
    Odrv4 I__608 (
            .O(N__3896),
            .I(\buart.Z_rx.startbit ));
    LocalMux I__607 (
            .O(N__3887),
            .I(\buart.Z_rx.startbit ));
    Odrv4 I__606 (
            .O(N__3884),
            .I(\buart.Z_rx.startbit ));
    LocalMux I__605 (
            .O(N__3875),
            .I(\buart.Z_rx.startbit ));
    LocalMux I__604 (
            .O(N__3872),
            .I(\buart.Z_rx.startbit ));
    LocalMux I__603 (
            .O(N__3869),
            .I(\buart.Z_rx.startbit ));
    CascadeMux I__602 (
            .O(N__3856),
            .I(N__3845));
    CascadeMux I__601 (
            .O(N__3855),
            .I(N__3841));
    InMux I__600 (
            .O(N__3854),
            .I(N__3838));
    InMux I__599 (
            .O(N__3853),
            .I(N__3835));
    InMux I__598 (
            .O(N__3852),
            .I(N__3832));
    InMux I__597 (
            .O(N__3851),
            .I(N__3827));
    InMux I__596 (
            .O(N__3850),
            .I(N__3827));
    InMux I__595 (
            .O(N__3849),
            .I(N__3822));
    InMux I__594 (
            .O(N__3848),
            .I(N__3822));
    InMux I__593 (
            .O(N__3845),
            .I(N__3815));
    InMux I__592 (
            .O(N__3844),
            .I(N__3815));
    InMux I__591 (
            .O(N__3841),
            .I(N__3815));
    LocalMux I__590 (
            .O(N__3838),
            .I(buart__rx_bitcount_2));
    LocalMux I__589 (
            .O(N__3835),
            .I(buart__rx_bitcount_2));
    LocalMux I__588 (
            .O(N__3832),
            .I(buart__rx_bitcount_2));
    LocalMux I__587 (
            .O(N__3827),
            .I(buart__rx_bitcount_2));
    LocalMux I__586 (
            .O(N__3822),
            .I(buart__rx_bitcount_2));
    LocalMux I__585 (
            .O(N__3815),
            .I(buart__rx_bitcount_2));
    InMux I__584 (
            .O(N__3802),
            .I(N__3799));
    LocalMux I__583 (
            .O(N__3799),
            .I(\Glue_Lab2.g0_8_2 ));
    InMux I__582 (
            .O(N__3796),
            .I(N__3793));
    LocalMux I__581 (
            .O(N__3793),
            .I(\Glue_Lab2.de0.un2_de_hexplusZ0Z_2 ));
    CascadeMux I__580 (
            .O(N__3790),
            .I(\Lab_UT.S_0_s_c2_1_cascade_ ));
    InMux I__579 (
            .O(N__3787),
            .I(N__3784));
    LocalMux I__578 (
            .O(N__3784),
            .I(\Lab_UT.S_0_s_ac0_5_0_2 ));
    InMux I__577 (
            .O(N__3781),
            .I(N__3778));
    LocalMux I__576 (
            .O(N__3778),
            .I(N__3775));
    Odrv4 I__575 (
            .O(N__3775),
            .I(Lab_UT_g1_1));
    InMux I__574 (
            .O(N__3772),
            .I(\buart.Z_rx.bitcount_cry_0 ));
    InMux I__573 (
            .O(N__3769),
            .I(\buart.Z_rx.bitcount_cry_1 ));
    InMux I__572 (
            .O(N__3766),
            .I(\buart.Z_rx.bitcount_cry_2 ));
    InMux I__571 (
            .O(N__3763),
            .I(\buart.Z_rx.bitcount_cry_3 ));
    InMux I__570 (
            .O(N__3760),
            .I(N__3757));
    LocalMux I__569 (
            .O(N__3757),
            .I(\buart.Z_rx.bitcount_lm_4 ));
    InMux I__568 (
            .O(N__3754),
            .I(N__3751));
    LocalMux I__567 (
            .O(N__3751),
            .I(\buart.Z_rx.bitcount_cry_0_THRU_CO ));
    InMux I__566 (
            .O(N__3748),
            .I(N__3745));
    LocalMux I__565 (
            .O(N__3745),
            .I(\buart.Z_rx.bitcount_cry_2_THRU_CO ));
    CascadeMux I__564 (
            .O(N__3742),
            .I(\buart.Z_rx.bitcount_lm_3_cascade_ ));
    InMux I__563 (
            .O(N__3739),
            .I(N__3736));
    LocalMux I__562 (
            .O(N__3736),
            .I(N__3733));
    Span4Mux_v I__561 (
            .O(N__3733),
            .I(N__3730));
    Odrv4 I__560 (
            .O(N__3730),
            .I(\Lab_UT.S_m_bm_N_5LZ0Z7 ));
    InMux I__559 (
            .O(N__3727),
            .I(N__3721));
    InMux I__558 (
            .O(N__3726),
            .I(N__3718));
    InMux I__557 (
            .O(N__3725),
            .I(N__3713));
    InMux I__556 (
            .O(N__3724),
            .I(N__3713));
    LocalMux I__555 (
            .O(N__3721),
            .I(Gl_r1_2_rep1));
    LocalMux I__554 (
            .O(N__3718),
            .I(Gl_r1_2_rep1));
    LocalMux I__553 (
            .O(N__3713),
            .I(Gl_r1_2_rep1));
    CascadeMux I__552 (
            .O(N__3706),
            .I(N__3700));
    CascadeMux I__551 (
            .O(N__3705),
            .I(N__3697));
    InMux I__550 (
            .O(N__3704),
            .I(N__3690));
    InMux I__549 (
            .O(N__3703),
            .I(N__3690));
    InMux I__548 (
            .O(N__3700),
            .I(N__3690));
    InMux I__547 (
            .O(N__3697),
            .I(N__3687));
    LocalMux I__546 (
            .O(N__3690),
            .I(N__3684));
    LocalMux I__545 (
            .O(N__3687),
            .I(Gl_r2_2_rep1));
    Odrv4 I__544 (
            .O(N__3684),
            .I(Gl_r2_2_rep1));
    InMux I__543 (
            .O(N__3679),
            .I(N__3676));
    LocalMux I__542 (
            .O(N__3676),
            .I(\Lab_UT.g0_4Z0Z_0 ));
    CEMux I__541 (
            .O(N__3673),
            .I(N__3669));
    CEMux I__540 (
            .O(N__3672),
            .I(N__3665));
    LocalMux I__539 (
            .O(N__3669),
            .I(N__3662));
    CEMux I__538 (
            .O(N__3668),
            .I(N__3659));
    LocalMux I__537 (
            .O(N__3665),
            .I(N__3656));
    Span4Mux_h I__536 (
            .O(N__3662),
            .I(N__3653));
    LocalMux I__535 (
            .O(N__3659),
            .I(N__3650));
    Span4Mux_v I__534 (
            .O(N__3656),
            .I(N__3647));
    Span4Mux_h I__533 (
            .O(N__3653),
            .I(N__3642));
    Span4Mux_h I__532 (
            .O(N__3650),
            .I(N__3642));
    Odrv4 I__531 (
            .O(N__3647),
            .I(\Glue_Lab2.Gl_r17_0_i ));
    Odrv4 I__530 (
            .O(N__3642),
            .I(\Glue_Lab2.Gl_r17_0_i ));
    InMux I__529 (
            .O(N__3637),
            .I(N__3634));
    LocalMux I__528 (
            .O(N__3634),
            .I(N__3631));
    Odrv4 I__527 (
            .O(N__3631),
            .I(\Lab_UT.g0_1_0_0 ));
    CEMux I__526 (
            .O(N__3628),
            .I(N__3624));
    CEMux I__525 (
            .O(N__3627),
            .I(N__3621));
    LocalMux I__524 (
            .O(N__3624),
            .I(\Glue_Lab2.Gl_r27_0_i ));
    LocalMux I__523 (
            .O(N__3621),
            .I(\Glue_Lab2.Gl_r27_0_i ));
    InMux I__522 (
            .O(N__3616),
            .I(N__3613));
    LocalMux I__521 (
            .O(N__3613),
            .I(\Lab_UT.g0_4_0_0 ));
    InMux I__520 (
            .O(N__3610),
            .I(N__3607));
    LocalMux I__519 (
            .O(N__3607),
            .I(\Lab_UT.S_1_ac0_1_0Z0Z_0 ));
    CascadeMux I__518 (
            .O(N__3604),
            .I(\Lab_UT.S_1_axbZ0Z1_cascade_ ));
    InMux I__517 (
            .O(N__3601),
            .I(N__3598));
    LocalMux I__516 (
            .O(N__3598),
            .I(\Lab_UT.g1Z0Z_0 ));
    CascadeMux I__515 (
            .O(N__3595),
            .I(\Lab_UT.S_0_s_c2_0_cascade_ ));
    InMux I__514 (
            .O(N__3592),
            .I(N__3589));
    LocalMux I__513 (
            .O(N__3589),
            .I(\Lab_UT.S_0_s_ac0_5_0_1 ));
    InMux I__512 (
            .O(N__3586),
            .I(N__3583));
    LocalMux I__511 (
            .O(N__3583),
            .I(\Lab_UT.gZ0Z1 ));
    CascadeMux I__510 (
            .O(N__3580),
            .I(N__3576));
    CascadeMux I__509 (
            .O(N__3579),
            .I(N__3573));
    InMux I__508 (
            .O(N__3576),
            .I(N__3567));
    InMux I__507 (
            .O(N__3573),
            .I(N__3567));
    InMux I__506 (
            .O(N__3572),
            .I(N__3564));
    LocalMux I__505 (
            .O(N__3567),
            .I(Glue_Lab2_Gl_r2_fast_0));
    LocalMux I__504 (
            .O(N__3564),
            .I(Glue_Lab2_Gl_r2_fast_0));
    InMux I__503 (
            .O(N__3559),
            .I(N__3552));
    InMux I__502 (
            .O(N__3558),
            .I(N__3552));
    CascadeMux I__501 (
            .O(N__3557),
            .I(N__3549));
    LocalMux I__500 (
            .O(N__3552),
            .I(N__3546));
    InMux I__499 (
            .O(N__3549),
            .I(N__3543));
    Odrv4 I__498 (
            .O(N__3546),
            .I(Glue_Lab2_Gl_r1_fast_0));
    LocalMux I__497 (
            .O(N__3543),
            .I(Glue_Lab2_Gl_r1_fast_0));
    CascadeMux I__496 (
            .O(N__3538),
            .I(\Glue_Lab2.gl_fsm.N_14_cascade_ ));
    InMux I__495 (
            .O(N__3535),
            .I(N__3528));
    InMux I__494 (
            .O(N__3534),
            .I(N__3528));
    CascadeMux I__493 (
            .O(N__3533),
            .I(N__3523));
    LocalMux I__492 (
            .O(N__3528),
            .I(N__3519));
    InMux I__491 (
            .O(N__3527),
            .I(N__3516));
    InMux I__490 (
            .O(N__3526),
            .I(N__3513));
    InMux I__489 (
            .O(N__3523),
            .I(N__3508));
    InMux I__488 (
            .O(N__3522),
            .I(N__3508));
    Span4Mux_s2_v I__487 (
            .O(N__3519),
            .I(N__3503));
    LocalMux I__486 (
            .O(N__3516),
            .I(N__3503));
    LocalMux I__485 (
            .O(N__3513),
            .I(Glue_Lab2_gl_fsm_state_0));
    LocalMux I__484 (
            .O(N__3508),
            .I(Glue_Lab2_gl_fsm_state_0));
    Odrv4 I__483 (
            .O(N__3503),
            .I(Glue_Lab2_gl_fsm_state_0));
    InMux I__482 (
            .O(N__3496),
            .I(N__3493));
    LocalMux I__481 (
            .O(N__3493),
            .I(\Lab_UT.C_out41_0 ));
    CascadeMux I__480 (
            .O(N__3490),
            .I(led_c_0_4_cascade_));
    CascadeMux I__479 (
            .O(N__3487),
            .I(N__3484));
    InMux I__478 (
            .O(N__3484),
            .I(N__3481));
    LocalMux I__477 (
            .O(N__3481),
            .I(N__3478));
    Odrv4 I__476 (
            .O(N__3478),
            .I(Gl_tx_data_6));
    InMux I__475 (
            .O(N__3475),
            .I(N__3472));
    LocalMux I__474 (
            .O(N__3472),
            .I(\Lab_UT.S_m_bm_N_2LZ0Z1 ));
    IoInMux I__473 (
            .O(N__3469),
            .I(N__3466));
    LocalMux I__472 (
            .O(N__3466),
            .I(N__3463));
    Span4Mux_s3_h I__471 (
            .O(N__3463),
            .I(N__3459));
    InMux I__470 (
            .O(N__3462),
            .I(N__3456));
    Odrv4 I__469 (
            .O(N__3459),
            .I(led_c_0));
    LocalMux I__468 (
            .O(N__3456),
            .I(led_c_0));
    CascadeMux I__467 (
            .O(N__3451),
            .I(bu_rx_data_rdy_cascade_));
    InMux I__466 (
            .O(N__3448),
            .I(N__3440));
    InMux I__465 (
            .O(N__3447),
            .I(N__3437));
    InMux I__464 (
            .O(N__3446),
            .I(N__3434));
    InMux I__463 (
            .O(N__3445),
            .I(N__3427));
    InMux I__462 (
            .O(N__3444),
            .I(N__3427));
    InMux I__461 (
            .O(N__3443),
            .I(N__3427));
    LocalMux I__460 (
            .O(N__3440),
            .I(N__3424));
    LocalMux I__459 (
            .O(N__3437),
            .I(N__3421));
    LocalMux I__458 (
            .O(N__3434),
            .I(\Glue_Lab2.i_rst_char_detected ));
    LocalMux I__457 (
            .O(N__3427),
            .I(\Glue_Lab2.i_rst_char_detected ));
    Odrv4 I__456 (
            .O(N__3424),
            .I(\Glue_Lab2.i_rst_char_detected ));
    Odrv4 I__455 (
            .O(N__3421),
            .I(\Glue_Lab2.i_rst_char_detected ));
    CascadeMux I__454 (
            .O(N__3412),
            .I(N__3409));
    InMux I__453 (
            .O(N__3409),
            .I(N__3404));
    InMux I__452 (
            .O(N__3408),
            .I(N__3401));
    InMux I__451 (
            .O(N__3407),
            .I(N__3398));
    LocalMux I__450 (
            .O(N__3404),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    LocalMux I__449 (
            .O(N__3401),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    LocalMux I__448 (
            .O(N__3398),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    CascadeMux I__447 (
            .O(N__3391),
            .I(N__3387));
    InMux I__446 (
            .O(N__3390),
            .I(N__3384));
    InMux I__445 (
            .O(N__3387),
            .I(N__3381));
    LocalMux I__444 (
            .O(N__3384),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ));
    LocalMux I__443 (
            .O(N__3381),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ));
    InMux I__442 (
            .O(N__3376),
            .I(N__3370));
    InMux I__441 (
            .O(N__3375),
            .I(N__3367));
    InMux I__440 (
            .O(N__3374),
            .I(N__3362));
    InMux I__439 (
            .O(N__3373),
            .I(N__3362));
    LocalMux I__438 (
            .O(N__3370),
            .I(N__3359));
    LocalMux I__437 (
            .O(N__3367),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ));
    LocalMux I__436 (
            .O(N__3362),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ));
    Odrv4 I__435 (
            .O(N__3359),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ));
    InMux I__434 (
            .O(N__3352),
            .I(N__3349));
    LocalMux I__433 (
            .O(N__3349),
            .I(N__3346));
    Odrv4 I__432 (
            .O(N__3346),
            .I(\buart.Z_rx.un1_sample_0 ));
    CascadeMux I__431 (
            .O(N__3343),
            .I(\buart.Z_rx.ser_clk_2_0_cascade_ ));
    CascadeMux I__430 (
            .O(N__3340),
            .I(\Glue_Lab2.de0.un2_de_hexplus_3_xZ0Z0_cascade_ ));
    CascadeMux I__429 (
            .O(N__3337),
            .I(\Glue_Lab2.de0.un2_de_hexplus_3_cascade_ ));
    CascadeMux I__428 (
            .O(N__3334),
            .I(\Glue_Lab2.is_hexplus_cascade_ ));
    InMux I__427 (
            .O(N__3331),
            .I(N__3328));
    LocalMux I__426 (
            .O(N__3328),
            .I(N__3325));
    Odrv4 I__425 (
            .O(N__3325),
            .I(Gl_tx_data_4));
    InMux I__424 (
            .O(N__3322),
            .I(N__3312));
    InMux I__423 (
            .O(N__3321),
            .I(N__3312));
    InMux I__422 (
            .O(N__3320),
            .I(N__3307));
    InMux I__421 (
            .O(N__3319),
            .I(N__3307));
    InMux I__420 (
            .O(N__3318),
            .I(N__3304));
    InMux I__419 (
            .O(N__3317),
            .I(N__3301));
    LocalMux I__418 (
            .O(N__3312),
            .I(\buart.Z_rx.ser_clk_2 ));
    LocalMux I__417 (
            .O(N__3307),
            .I(\buart.Z_rx.ser_clk_2 ));
    LocalMux I__416 (
            .O(N__3304),
            .I(\buart.Z_rx.ser_clk_2 ));
    LocalMux I__415 (
            .O(N__3301),
            .I(\buart.Z_rx.ser_clk_2 ));
    CascadeMux I__414 (
            .O(N__3292),
            .I(N__3288));
    CascadeMux I__413 (
            .O(N__3291),
            .I(N__3285));
    InMux I__412 (
            .O(N__3288),
            .I(N__3280));
    InMux I__411 (
            .O(N__3285),
            .I(N__3277));
    InMux I__410 (
            .O(N__3284),
            .I(N__3274));
    InMux I__409 (
            .O(N__3283),
            .I(N__3271));
    LocalMux I__408 (
            .O(N__3280),
            .I(N__3268));
    LocalMux I__407 (
            .O(N__3277),
            .I(\buart.Z_rx.ser_clk_2_0 ));
    LocalMux I__406 (
            .O(N__3274),
            .I(\buart.Z_rx.ser_clk_2_0 ));
    LocalMux I__405 (
            .O(N__3271),
            .I(\buart.Z_rx.ser_clk_2_0 ));
    Odrv4 I__404 (
            .O(N__3268),
            .I(\buart.Z_rx.ser_clk_2_0 ));
    CascadeMux I__403 (
            .O(N__3259),
            .I(N__3255));
    CascadeMux I__402 (
            .O(N__3258),
            .I(N__3250));
    InMux I__401 (
            .O(N__3255),
            .I(N__3246));
    InMux I__400 (
            .O(N__3254),
            .I(N__3241));
    InMux I__399 (
            .O(N__3253),
            .I(N__3241));
    InMux I__398 (
            .O(N__3250),
            .I(N__3236));
    InMux I__397 (
            .O(N__3249),
            .I(N__3236));
    LocalMux I__396 (
            .O(N__3246),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    LocalMux I__395 (
            .O(N__3241),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    LocalMux I__394 (
            .O(N__3236),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    CascadeMux I__393 (
            .O(N__3229),
            .I(N__3226));
    InMux I__392 (
            .O(N__3226),
            .I(N__3223));
    LocalMux I__391 (
            .O(N__3223),
            .I(\Glue_Lab2.de0.g0_5_0 ));
    InMux I__390 (
            .O(N__3220),
            .I(N__3217));
    LocalMux I__389 (
            .O(N__3217),
            .I(N__3214));
    Span4Mux_h I__388 (
            .O(N__3214),
            .I(N__3208));
    InMux I__387 (
            .O(N__3213),
            .I(N__3205));
    InMux I__386 (
            .O(N__3212),
            .I(N__3200));
    InMux I__385 (
            .O(N__3211),
            .I(N__3200));
    Odrv4 I__384 (
            .O(N__3208),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__383 (
            .O(N__3205),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__382 (
            .O(N__3200),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    InMux I__381 (
            .O(N__3193),
            .I(N__3188));
    InMux I__380 (
            .O(N__3192),
            .I(N__3185));
    InMux I__379 (
            .O(N__3191),
            .I(N__3182));
    LocalMux I__378 (
            .O(N__3188),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ));
    LocalMux I__377 (
            .O(N__3185),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ));
    LocalMux I__376 (
            .O(N__3182),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ));
    CascadeMux I__375 (
            .O(N__3175),
            .I(\Glue_Lab2.de0.g0_5_2_cascade_ ));
    CascadeMux I__374 (
            .O(N__3172),
            .I(\Glue_Lab2.g0_9_2_cascade_ ));
    InMux I__373 (
            .O(N__3169),
            .I(N__3166));
    LocalMux I__372 (
            .O(N__3166),
            .I(N__3163));
    Odrv4 I__371 (
            .O(N__3163),
            .I(\Glue_Lab2.g0_7_2 ));
    InMux I__370 (
            .O(N__3160),
            .I(N__3157));
    LocalMux I__369 (
            .O(N__3157),
            .I(\Glue_Lab2.reset_counte_0_3 ));
    CascadeMux I__368 (
            .O(N__3154),
            .I(\buart.Z_rx.bitcount_RNIMK771_0Z0Z_4_cascade_ ));
    CascadeMux I__367 (
            .O(N__3151),
            .I(\Glue_Lab2.g0_9_0_cascade_ ));
    InMux I__366 (
            .O(N__3148),
            .I(N__3145));
    LocalMux I__365 (
            .O(N__3145),
            .I(\Glue_Lab2.reset_counte_0_1 ));
    InMux I__364 (
            .O(N__3142),
            .I(N__3139));
    LocalMux I__363 (
            .O(N__3139),
            .I(\Glue_Lab2.g0_7_0 ));
    CascadeMux I__362 (
            .O(N__3136),
            .I(\buart.Z_rx.bitcountlde_0_cascade_ ));
    IoInMux I__361 (
            .O(N__3133),
            .I(N__3130));
    LocalMux I__360 (
            .O(N__3130),
            .I(N__3126));
    CascadeMux I__359 (
            .O(N__3129),
            .I(N__3123));
    Span4Mux_s3_v I__358 (
            .O(N__3126),
            .I(N__3120));
    InMux I__357 (
            .O(N__3123),
            .I(N__3116));
    Span4Mux_v I__356 (
            .O(N__3120),
            .I(N__3113));
    InMux I__355 (
            .O(N__3119),
            .I(N__3110));
    LocalMux I__354 (
            .O(N__3116),
            .I(N__3107));
    Span4Mux_h I__353 (
            .O(N__3113),
            .I(N__3104));
    LocalMux I__352 (
            .O(N__3110),
            .I(N__3099));
    Span4Mux_h I__351 (
            .O(N__3107),
            .I(N__3099));
    Odrv4 I__350 (
            .O(N__3104),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__349 (
            .O(N__3099),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__348 (
            .O(N__3094),
            .I(\buart.Z_rx.N_29_0_i_cascade_ ));
    InMux I__347 (
            .O(N__3091),
            .I(N__3088));
    LocalMux I__346 (
            .O(N__3088),
            .I(\buart.Z_rx.bitcount_lm_0 ));
    CascadeMux I__345 (
            .O(N__3085),
            .I(N__3082));
    InMux I__344 (
            .O(N__3082),
            .I(N__3079));
    LocalMux I__343 (
            .O(N__3079),
            .I(N__3076));
    Odrv12 I__342 (
            .O(N__3076),
            .I(\Lab_UT.S_m_bm_N_6LZ0Z10 ));
    CascadeMux I__341 (
            .O(N__3073),
            .I(\Lab_UT.g0_0_a3Z0Z_0_cascade_ ));
    InMux I__340 (
            .O(N__3070),
            .I(N__3067));
    LocalMux I__339 (
            .O(N__3067),
            .I(\Lab_UT.g0_1Z0Z_0 ));
    InMux I__338 (
            .O(N__3064),
            .I(N__3061));
    LocalMux I__337 (
            .O(N__3061),
            .I(\Lab_UT.N_6 ));
    CascadeMux I__336 (
            .O(N__3058),
            .I(\Lab_UT.S_0_s_axbZ0Z3_cascade_ ));
    InMux I__335 (
            .O(N__3055),
            .I(N__3052));
    LocalMux I__334 (
            .O(N__3052),
            .I(N__3049));
    Odrv4 I__333 (
            .O(N__3049),
            .I(\Lab_UT.S_m_amZ0Z_3 ));
    InMux I__332 (
            .O(N__3046),
            .I(N__3043));
    LocalMux I__331 (
            .O(N__3043),
            .I(N__3040));
    Odrv12 I__330 (
            .O(N__3040),
            .I(\Lab_UT.g1_0_0 ));
    CascadeMux I__329 (
            .O(N__3037),
            .I(\Lab_UT.S_m_bmZ0Z_3_cascade_ ));
    IoInMux I__328 (
            .O(N__3034),
            .I(N__3031));
    LocalMux I__327 (
            .O(N__3031),
            .I(N__3028));
    IoSpan4Mux I__326 (
            .O(N__3028),
            .I(N__3025));
    Span4Mux_s3_h I__325 (
            .O(N__3025),
            .I(N__3022));
    Odrv4 I__324 (
            .O(N__3022),
            .I(led_c_3));
    CascadeMux I__323 (
            .O(N__3019),
            .I(led_c_3_cascade_));
    InMux I__322 (
            .O(N__3016),
            .I(N__3013));
    LocalMux I__321 (
            .O(N__3013),
            .I(N__3010));
    Odrv4 I__320 (
            .O(N__3010),
            .I(Gl_tx_data_3));
    InMux I__319 (
            .O(N__3007),
            .I(N__3004));
    LocalMux I__318 (
            .O(N__3004),
            .I(\Lab_UT.S_m_bm_N_3LZ0Z3 ));
    CascadeMux I__317 (
            .O(N__3001),
            .I(\Lab_UT.g0_0_a3_0Z0Z_0_cascade_ ));
    CascadeMux I__316 (
            .O(N__2998),
            .I(Lab_UT_C_out41_1_cascade_));
    InMux I__315 (
            .O(N__2995),
            .I(N__2992));
    LocalMux I__314 (
            .O(N__2992),
            .I(N__2989));
    Odrv12 I__313 (
            .O(N__2989),
            .I(Gl_tx_data_5));
    InMux I__312 (
            .O(N__2986),
            .I(N__2983));
    LocalMux I__311 (
            .O(N__2983),
            .I(\Lab_UT.N_6_0 ));
    InMux I__310 (
            .O(N__2980),
            .I(N__2977));
    LocalMux I__309 (
            .O(N__2977),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_ac0_7 ));
    CascadeMux I__308 (
            .O(N__2974),
            .I(\buart.Z_rx.ser_clk_2_cascade_ ));
    InMux I__307 (
            .O(N__2971),
            .I(N__2967));
    InMux I__306 (
            .O(N__2970),
            .I(N__2964));
    LocalMux I__305 (
            .O(N__2967),
            .I(\Glue_Lab2.reset_countZ0Z_0 ));
    LocalMux I__304 (
            .O(N__2964),
            .I(\Glue_Lab2.reset_countZ0Z_0 ));
    InMux I__303 (
            .O(N__2959),
            .I(N__2956));
    LocalMux I__302 (
            .O(N__2956),
            .I(\buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_4 ));
    InMux I__301 (
            .O(N__2953),
            .I(N__2950));
    LocalMux I__300 (
            .O(N__2950),
            .I(\Lab_UT.sDelay.delayRegZ0Z_0 ));
    InMux I__299 (
            .O(N__2947),
            .I(N__2944));
    LocalMux I__298 (
            .O(N__2944),
            .I(N__2941));
    Odrv4 I__297 (
            .O(N__2941),
            .I(Gl_tx_data_0));
    InMux I__296 (
            .O(N__2938),
            .I(N__2935));
    LocalMux I__295 (
            .O(N__2935),
            .I(\buart.Z_tx.shifterZ0Z_2 ));
    InMux I__294 (
            .O(N__2932),
            .I(N__2929));
    LocalMux I__293 (
            .O(N__2929),
            .I(\buart.Z_tx.shifterZ0Z_3 ));
    InMux I__292 (
            .O(N__2926),
            .I(N__2923));
    LocalMux I__291 (
            .O(N__2923),
            .I(\buart.Z_tx.shifterZ0Z_4 ));
    InMux I__290 (
            .O(N__2920),
            .I(N__2917));
    LocalMux I__289 (
            .O(N__2917),
            .I(\buart.Z_tx.shifterZ0Z_5 ));
    InMux I__288 (
            .O(N__2914),
            .I(N__2911));
    LocalMux I__287 (
            .O(N__2911),
            .I(\buart.Z_tx.shifterZ0Z_7 ));
    InMux I__286 (
            .O(N__2908),
            .I(N__2905));
    LocalMux I__285 (
            .O(N__2905),
            .I(\buart.Z_tx.shifterZ0Z_6 ));
    InMux I__284 (
            .O(N__2902),
            .I(N__2899));
    LocalMux I__283 (
            .O(N__2899),
            .I(\Glue_Lab2.reset_count_cry_2_THRU_CO ));
    CascadeMux I__282 (
            .O(N__2896),
            .I(N__2893));
    InMux I__281 (
            .O(N__2893),
            .I(N__2889));
    InMux I__280 (
            .O(N__2892),
            .I(N__2886));
    LocalMux I__279 (
            .O(N__2889),
            .I(\Glue_Lab2.reset_countZ0Z_3 ));
    LocalMux I__278 (
            .O(N__2886),
            .I(\Glue_Lab2.reset_countZ0Z_3 ));
    CascadeMux I__277 (
            .O(N__2881),
            .I(N__2878));
    InMux I__276 (
            .O(N__2878),
            .I(N__2875));
    LocalMux I__275 (
            .O(N__2875),
            .I(\Glue_Lab2.reset_count_cry_0_THRU_CO ));
    InMux I__274 (
            .O(N__2872),
            .I(N__2868));
    InMux I__273 (
            .O(N__2871),
            .I(N__2865));
    LocalMux I__272 (
            .O(N__2868),
            .I(\Glue_Lab2.reset_countZ0Z_1 ));
    LocalMux I__271 (
            .O(N__2865),
            .I(\Glue_Lab2.reset_countZ0Z_1 ));
    CascadeMux I__270 (
            .O(N__2860),
            .I(\buart.Z_rx.Z_baudgen.counter_0_1_5_cascade_ ));
    InMux I__269 (
            .O(N__2857),
            .I(\Glue_Lab2.reset_count_cry_1 ));
    InMux I__268 (
            .O(N__2854),
            .I(\Glue_Lab2.reset_count_cry_2 ));
    InMux I__267 (
            .O(N__2851),
            .I(\Glue_Lab2.reset_count_cry_3 ));
    InMux I__266 (
            .O(N__2848),
            .I(N__2845));
    LocalMux I__265 (
            .O(N__2845),
            .I(N__2842));
    Odrv4 I__264 (
            .O(N__2842),
            .I(\Glue_Lab2.reset_count_cry_1_THRU_CO ));
    CascadeMux I__263 (
            .O(N__2839),
            .I(N__2835));
    CascadeMux I__262 (
            .O(N__2838),
            .I(N__2832));
    InMux I__261 (
            .O(N__2835),
            .I(N__2829));
    InMux I__260 (
            .O(N__2832),
            .I(N__2826));
    LocalMux I__259 (
            .O(N__2829),
            .I(N__2823));
    LocalMux I__258 (
            .O(N__2826),
            .I(\Glue_Lab2.reset_countZ0Z_2 ));
    Odrv4 I__257 (
            .O(N__2823),
            .I(\Glue_Lab2.reset_countZ0Z_2 ));
    InMux I__256 (
            .O(N__2818),
            .I(N__2815));
    LocalMux I__255 (
            .O(N__2815),
            .I(\buart.Z_tx.shifterZ0Z_1 ));
    InMux I__254 (
            .O(N__2812),
            .I(N__2809));
    LocalMux I__253 (
            .O(N__2809),
            .I(\buart.Z_tx.shifterZ0Z_0 ));
    IoInMux I__252 (
            .O(N__2806),
            .I(N__2803));
    LocalMux I__251 (
            .O(N__2803),
            .I(N__2800));
    IoSpan4Mux I__250 (
            .O(N__2800),
            .I(N__2797));
    Odrv4 I__249 (
            .O(N__2797),
            .I(clk_in_c));
    IoInMux I__248 (
            .O(N__2794),
            .I(N__2791));
    LocalMux I__247 (
            .O(N__2791),
            .I(N__2788));
    Span4Mux_s1_h I__246 (
            .O(N__2788),
            .I(N__2785));
    Span4Mux_h I__245 (
            .O(N__2785),
            .I(N__2782));
    Sp12to4 I__244 (
            .O(N__2782),
            .I(N__2779));
    Odrv12 I__243 (
            .O(N__2779),
            .I(clk));
    InMux I__242 (
            .O(N__2776),
            .I(N__2773));
    LocalMux I__241 (
            .O(N__2773),
            .I(N__2770));
    Span4Mux_h I__240 (
            .O(N__2770),
            .I(N__2767));
    IoSpan4Mux I__239 (
            .O(N__2767),
            .I(N__2764));
    Odrv4 I__238 (
            .O(N__2764),
            .I(uart_RXD));
    IoInMux I__237 (
            .O(N__2761),
            .I(N__2758));
    LocalMux I__236 (
            .O(N__2758),
            .I(N__2755));
    IoSpan4Mux I__235 (
            .O(N__2755),
            .I(N__2752));
    Span4Mux_s3_h I__234 (
            .O(N__2752),
            .I(N__2749));
    Odrv4 I__233 (
            .O(N__2749),
            .I(o_serial_data_c));
    InMux I__232 (
            .O(N__2746),
            .I(\Glue_Lab2.reset_count_cry_0 ));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_9_0_));
    defparam IN_MUX_bfv_6_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_11_0_));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB clk_derived_clock_RNI7BQ7 (
            .USERSIGNALTOGLOBALBUFFER(N__2794),
            .GLOBALBUFFEROUTPUT(clk_g));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \buart.Z_rx.hh_1_LC_5_10_1 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_1_LC_5_10_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.hh_1_LC_5_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.hh_1_LC_5_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4059),
            .lcout(\buart.Z_rx.hhZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6163),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.hh_0_LC_5_10_6 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_0_LC_5_10_6 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.hh_0_LC_5_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.hh_0_LC_5_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2776),
            .lcout(\buart.Z_rx.hhZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6163),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.uart_tx_LC_6_10_6 .C_ON=1'b0;
    defparam \buart.Z_tx.uart_tx_LC_6_10_6 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.uart_tx_LC_6_10_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \buart.Z_tx.uart_tx_LC_6_10_6  (
            .in0(_gnd_net_),
            .in1(N__2812),
            .in2(_gnd_net_),
            .in3(N__6796),
            .lcout(o_serial_data_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6165),
            .ce(N__6711),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.reset_count_cry_c_0_LC_6_11_0 .C_ON=1'b1;
    defparam \Glue_Lab2.reset_count_cry_c_0_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.reset_count_cry_c_0_LC_6_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \Glue_Lab2.reset_count_cry_c_0_LC_6_11_0  (
            .in0(_gnd_net_),
            .in1(N__2970),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_11_0_),
            .carryout(\Glue_Lab2.reset_count_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.reset_count_cry_0_THRU_LUT4_0_LC_6_11_1 .C_ON=1'b1;
    defparam \Glue_Lab2.reset_count_cry_0_THRU_LUT4_0_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.reset_count_cry_0_THRU_LUT4_0_LC_6_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Glue_Lab2.reset_count_cry_0_THRU_LUT4_0_LC_6_11_1  (
            .in0(_gnd_net_),
            .in1(N__2871),
            .in2(_gnd_net_),
            .in3(N__2746),
            .lcout(\Glue_Lab2.reset_count_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\Glue_Lab2.reset_count_cry_0 ),
            .carryout(\Glue_Lab2.reset_count_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.reset_count_cry_1_THRU_LUT4_0_LC_6_11_2 .C_ON=1'b1;
    defparam \Glue_Lab2.reset_count_cry_1_THRU_LUT4_0_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.reset_count_cry_1_THRU_LUT4_0_LC_6_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Glue_Lab2.reset_count_cry_1_THRU_LUT4_0_LC_6_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2839),
            .in3(N__2857),
            .lcout(\Glue_Lab2.reset_count_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\Glue_Lab2.reset_count_cry_1 ),
            .carryout(\Glue_Lab2.reset_count_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.reset_count_cry_2_THRU_LUT4_0_LC_6_11_3 .C_ON=1'b1;
    defparam \Glue_Lab2.reset_count_cry_2_THRU_LUT4_0_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.reset_count_cry_2_THRU_LUT4_0_LC_6_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Glue_Lab2.reset_count_cry_2_THRU_LUT4_0_LC_6_11_3  (
            .in0(_gnd_net_),
            .in1(N__2892),
            .in2(_gnd_net_),
            .in3(N__2854),
            .lcout(\Glue_Lab2.reset_count_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\Glue_Lab2.reset_count_cry_2 ),
            .carryout(\Glue_Lab2.reset_count_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.reset_count_4_LC_6_11_4 .C_ON=1'b0;
    defparam \Glue_Lab2.reset_count_4_LC_6_11_4 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.reset_count_4_LC_6_11_4 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \Glue_Lab2.reset_count_4_LC_6_11_4  (
            .in0(N__3447),
            .in1(N__5292),
            .in2(_gnd_net_),
            .in3(N__2851),
            .lcout(\Glue_Lab2.reset_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6166),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_6_11_5 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_6_11_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_6_11_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_0_LC_6_11_5  (
            .in0(_gnd_net_),
            .in1(N__3213),
            .in2(_gnd_net_),
            .in3(N__3946),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6166),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_7_8_6.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_7_8_6.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_7_8_6.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_7_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.reset_count_2_LC_7_9_1 .C_ON=1'b0;
    defparam \Glue_Lab2.reset_count_2_LC_7_9_1 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.reset_count_2_LC_7_9_1 .LUT_INIT=16'b1100000011010010;
    LogicCell40 \Glue_Lab2.reset_count_2_LC_7_9_1  (
            .in0(N__2848),
            .in1(N__3148),
            .in2(N__2838),
            .in3(N__3448),
            .lcout(\Glue_Lab2.reset_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6164),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_1_LC_7_10_0 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_1_LC_7_10_0 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.shifter_1_LC_7_10_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_1_LC_7_10_0  (
            .in0(N__6789),
            .in1(N__2938),
            .in2(_gnd_net_),
            .in3(N__2947),
            .lcout(\buart.Z_tx.shifterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6167),
            .ce(N__6715),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_0_LC_7_10_1 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_0_LC_7_10_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.shifter_0_LC_7_10_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \buart.Z_tx.shifter_0_LC_7_10_1  (
            .in0(_gnd_net_),
            .in1(N__6788),
            .in2(_gnd_net_),
            .in3(N__2818),
            .lcout(\buart.Z_tx.shifterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6167),
            .ce(N__6715),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_7_LC_7_10_2 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_7_LC_7_10_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.shifter_7_LC_7_10_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \buart.Z_tx.shifter_7_LC_7_10_2  (
            .in0(N__6795),
            .in1(_gnd_net_),
            .in2(N__3487),
            .in3(N__6727),
            .lcout(\buart.Z_tx.shifterZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6167),
            .ce(N__6715),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_2_LC_7_10_3 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_2_LC_7_10_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.shifter_2_LC_7_10_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \buart.Z_tx.shifter_2_LC_7_10_3  (
            .in0(N__2932),
            .in1(N__6790),
            .in2(_gnd_net_),
            .in3(N__4762),
            .lcout(\buart.Z_tx.shifterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6167),
            .ce(N__6715),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_3_LC_7_10_4 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_3_LC_7_10_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.shifter_3_LC_7_10_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_3_LC_7_10_4  (
            .in0(N__6791),
            .in1(N__2926),
            .in2(_gnd_net_),
            .in3(N__4249),
            .lcout(\buart.Z_tx.shifterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6167),
            .ce(N__6715),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_4_LC_7_10_5 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_4_LC_7_10_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.shifter_4_LC_7_10_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \buart.Z_tx.shifter_4_LC_7_10_5  (
            .in0(N__2920),
            .in1(N__6792),
            .in2(_gnd_net_),
            .in3(N__3016),
            .lcout(\buart.Z_tx.shifterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6167),
            .ce(N__6715),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_5_LC_7_10_6 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_5_LC_7_10_6 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.shifter_5_LC_7_10_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \buart.Z_tx.shifter_5_LC_7_10_6  (
            .in0(N__6793),
            .in1(N__3331),
            .in2(_gnd_net_),
            .in3(N__2908),
            .lcout(\buart.Z_tx.shifterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6167),
            .ce(N__6715),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_6_LC_7_10_7 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_6_LC_7_10_7 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.shifter_6_LC_7_10_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \buart.Z_tx.shifter_6_LC_7_10_7  (
            .in0(N__2914),
            .in1(N__6794),
            .in2(_gnd_net_),
            .in3(N__2995),
            .lcout(\buart.Z_tx.shifterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6167),
            .ce(N__6715),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.reset_count_3_LC_7_11_0 .C_ON=1'b0;
    defparam \Glue_Lab2.reset_count_3_LC_7_11_0 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.reset_count_3_LC_7_11_0 .LUT_INIT=16'b1111000000010100;
    LogicCell40 \Glue_Lab2.reset_count_3_LC_7_11_0  (
            .in0(N__3443),
            .in1(N__2902),
            .in2(N__2896),
            .in3(N__5248),
            .lcout(\Glue_Lab2.reset_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6168),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.reset_count_1_LC_7_11_1 .C_ON=1'b0;
    defparam \Glue_Lab2.reset_count_1_LC_7_11_1 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.reset_count_1_LC_7_11_1 .LUT_INIT=16'b1000100010011010;
    LogicCell40 \Glue_Lab2.reset_count_1_LC_7_11_1  (
            .in0(N__2872),
            .in1(N__5509),
            .in2(N__2881),
            .in3(N__3445),
            .lcout(\Glue_Lab2.reset_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6168),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNO_0_5_LC_7_11_2 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNO_0_5_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNO_0_5_LC_7_11_2 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNO_0_5_LC_7_11_2  (
            .in0(N__3212),
            .in1(N__3192),
            .in2(_gnd_net_),
            .in3(N__3283),
            .lcout(),
            .ltout(\buart.Z_rx.Z_baudgen.counter_0_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_7_11_3 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_7_11_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_7_11_3 .LUT_INIT=16'b0000000001100000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_5_LC_7_11_3  (
            .in0(N__3390),
            .in1(N__2980),
            .in2(N__2860),
            .in3(N__3945),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6168),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNO_1_5_LC_7_11_4 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNO_1_5_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNO_1_5_LC_7_11_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNO_1_5_LC_7_11_4  (
            .in0(N__3374),
            .in1(N__3254),
            .in2(N__3412),
            .in3(N__3318),
            .lcout(\buart.Z_rx.Z_baudgen.un5_counter_ac0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNIT3N1_1_LC_7_11_5 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNIT3N1_1_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNIT3N1_1_LC_7_11_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNIT3N1_1_LC_7_11_5  (
            .in0(_gnd_net_),
            .in1(N__3191),
            .in2(_gnd_net_),
            .in3(N__3211),
            .lcout(\buart.Z_rx.ser_clk_2 ),
            .ltout(\buart.Z_rx.ser_clk_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNO_0_4_LC_7_11_6 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNO_0_4_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNO_0_4_LC_7_11_6 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNO_0_4_LC_7_11_6  (
            .in0(N__3373),
            .in1(N__3408),
            .in2(N__2974),
            .in3(N__3253),
            .lcout(\buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.reset_count_0_LC_7_11_7 .C_ON=1'b0;
    defparam \Glue_Lab2.reset_count_0_LC_7_11_7 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.reset_count_0_LC_7_11_7 .LUT_INIT=16'b1000100010011010;
    LogicCell40 \Glue_Lab2.reset_count_0_LC_7_11_7  (
            .in0(N__2971),
            .in1(N__3160),
            .in2(N__3129),
            .in3(N__3444),
            .lcout(\Glue_Lab2.reset_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6168),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.sDelay.delayReg_1_LC_7_12_1 .C_ON=1'b0;
    defparam \Lab_UT.sDelay.delayReg_1_LC_7_12_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.sDelay.delayReg_1_LC_7_12_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \Lab_UT.sDelay.delayReg_1_LC_7_12_1  (
            .in0(N__2953),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6247),
            .lcout(\Lab_UT.sDelay.delayRegZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6170),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_7_12_2 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_7_12_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_7_12_2 .LUT_INIT=16'b0000010001000100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_4_LC_7_12_2  (
            .in0(N__3943),
            .in1(N__2959),
            .in2(N__3291),
            .in3(N__3321),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6170),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_7_12_3 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_7_12_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_7_12_3 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_3_LC_7_12_3  (
            .in0(N__3322),
            .in1(N__3375),
            .in2(N__3259),
            .in3(N__3944),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6170),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.sDelay.delayReg_0_LC_7_12_4 .C_ON=1'b0;
    defparam \Lab_UT.sDelay.delayReg_0_LC_7_12_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.sDelay.delayReg_0_LC_7_12_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.sDelay.delayReg_0_LC_7_12_4  (
            .in0(N__6246),
            .in1(N__4697),
            .in2(_gnd_net_),
            .in3(N__3526),
            .lcout(\Lab_UT.sDelay.delayRegZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6170),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_tx_data_0_LC_7_12_5 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_tx_data_0_LC_7_12_5 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.Gl_tx_data_0_LC_7_12_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Glue_Lab2.Gl_tx_data_0_LC_7_12_5  (
            .in0(N__3462),
            .in1(N__5382),
            .in2(_gnd_net_),
            .in3(N__5016),
            .lcout(Gl_tx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6170),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_rst_LC_7_12_7 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_rst_LC_7_12_7 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.Gl_rst_LC_7_12_7 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \Glue_Lab2.Gl_rst_LC_7_12_7  (
            .in0(N__5293),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3446),
            .lcout(Gl_rst),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6170),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.S_m_bm_3_LC_7_13_0 .C_ON=1'b0;
    defparam \Lab_UT.S_m_bm_3_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.S_m_bm_3_LC_7_13_0 .LUT_INIT=16'b1100110001100011;
    LogicCell40 \Lab_UT.S_m_bm_3_LC_7_13_0  (
            .in0(N__3739),
            .in1(N__3007),
            .in2(N__3085),
            .in3(N__3475),
            .lcout(),
            .ltout(\Lab_UT.S_m_bmZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.S_m_ns_3_LC_7_13_1 .C_ON=1'b0;
    defparam \Lab_UT.S_m_ns_3_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.S_m_ns_3_LC_7_13_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \Lab_UT.S_m_ns_3_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(N__3055),
            .in2(N__3037),
            .in3(N__5571),
            .lcout(led_c_3),
            .ltout(led_c_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_tx_data_3_LC_7_13_2 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_tx_data_3_LC_7_13_2 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.Gl_tx_data_3_LC_7_13_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \Glue_Lab2.Gl_tx_data_3_LC_7_13_2  (
            .in0(_gnd_net_),
            .in1(N__6614),
            .in2(N__3019),
            .in3(N__5017),
            .lcout(Gl_tx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6173),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.S_m_bm_N_3L3_LC_7_13_3 .C_ON=1'b0;
    defparam \Lab_UT.S_m_bm_N_3L3_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.S_m_bm_N_3L3_LC_7_13_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.S_m_bm_N_3L3_LC_7_13_3  (
            .in0(_gnd_net_),
            .in1(N__5651),
            .in2(_gnd_net_),
            .in3(N__5718),
            .lcout(\Lab_UT.S_m_bm_N_3LZ0Z3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.g0_0_a3_0_1_LC_7_13_4 .C_ON=1'b0;
    defparam \Lab_UT.g0_0_a3_0_1_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.g0_0_a3_0_1_LC_7_13_4 .LUT_INIT=16'b1010111100100011;
    LogicCell40 \Lab_UT.g0_0_a3_0_1_LC_7_13_4  (
            .in0(N__5720),
            .in1(N__5813),
            .in2(N__5661),
            .in3(N__5882),
            .lcout(),
            .ltout(\Lab_UT.g0_0_a3_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.g0_1_LC_7_13_5 .C_ON=1'b0;
    defparam \Lab_UT.g0_1_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.g0_1_LC_7_13_5 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \Lab_UT.g0_1_LC_7_13_5  (
            .in0(N__3637),
            .in1(N__3046),
            .in2(N__3001),
            .in3(N__2986),
            .lcout(),
            .ltout(Lab_UT_C_out41_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_tx_data_5_LC_7_13_6 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_tx_data_5_LC_7_13_6 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.Gl_tx_data_5_LC_7_13_6 .LUT_INIT=16'b1111111111010001;
    LogicCell40 \Glue_Lab2.Gl_tx_data_5_LC_7_13_6  (
            .in0(N__3781),
            .in1(N__5896),
            .in2(N__2998),
            .in3(N__5018),
            .lcout(Gl_tx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6173),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.g0_0_a3_LC_7_13_7 .C_ON=1'b0;
    defparam \Lab_UT.g0_0_a3_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.g0_0_a3_LC_7_13_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.g0_0_a3_LC_7_13_7  (
            .in0(_gnd_net_),
            .in1(N__5652),
            .in2(_gnd_net_),
            .in3(N__5719),
            .lcout(\Lab_UT.N_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_r1_1_LC_7_14_1 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_r1_1_LC_7_14_1 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.Gl_r1_1_LC_7_14_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Glue_Lab2.Gl_r1_1_LC_7_14_1  (
            .in0(N__6352),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6474),
            .lcout(Gl_r1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6178),
            .ce(N__3668),
            .sr(_gnd_net_));
    defparam \Lab_UT.g0_0_a3_0_0_LC_7_14_2 .C_ON=1'b0;
    defparam \Lab_UT.g0_0_a3_0_0_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.g0_0_a3_0_0_LC_7_14_2 .LUT_INIT=16'b1010111100100011;
    LogicCell40 \Lab_UT.g0_0_a3_0_0_LC_7_14_2  (
            .in0(N__5717),
            .in1(N__3704),
            .in2(N__5656),
            .in3(N__3725),
            .lcout(),
            .ltout(\Lab_UT.g0_0_a3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.g0_0_LC_7_14_3 .C_ON=1'b0;
    defparam \Lab_UT.g0_0_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.g0_0_LC_7_14_3 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \Lab_UT.g0_0_LC_7_14_3  (
            .in0(N__3601),
            .in1(N__3070),
            .in2(N__3073),
            .in3(N__3064),
            .lcout(\Lab_UT.C_out41_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.g0_1_0_LC_7_14_4 .C_ON=1'b0;
    defparam \Lab_UT.g0_1_0_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.g0_1_0_LC_7_14_4 .LUT_INIT=16'b0011000010111010;
    LogicCell40 \Lab_UT.g0_1_0_LC_7_14_4  (
            .in0(N__3726),
            .in1(N__4549),
            .in2(N__4414),
            .in3(N__3703),
            .lcout(\Lab_UT.g0_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.g0_0_a3_0_LC_7_14_5 .C_ON=1'b0;
    defparam \Lab_UT.g0_0_a3_0_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.g0_0_a3_0_LC_7_14_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.g0_0_a3_0_LC_7_14_5  (
            .in0(_gnd_net_),
            .in1(N__5642),
            .in2(_gnd_net_),
            .in3(N__5715),
            .lcout(\Lab_UT.N_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_r1_3_LC_7_14_6 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_r1_3_LC_7_14_6 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.Gl_r1_3_LC_7_14_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Glue_Lab2.Gl_r1_3_LC_7_14_6  (
            .in0(_gnd_net_),
            .in1(N__6353),
            .in2(_gnd_net_),
            .in3(N__6615),
            .lcout(Gl_r1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6178),
            .ce(N__3668),
            .sr(_gnd_net_));
    defparam \Lab_UT.g0_3_LC_7_14_7 .C_ON=1'b0;
    defparam \Lab_UT.g0_3_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.g0_3_LC_7_14_7 .LUT_INIT=16'b1110110010000000;
    LogicCell40 \Lab_UT.g0_3_LC_7_14_7  (
            .in0(N__3724),
            .in1(N__5641),
            .in2(N__3706),
            .in3(N__5716),
            .lcout(\Lab_UT.S_0_s_ac0_5_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.S_0_s_axb3_LC_7_15_0 .C_ON=1'b0;
    defparam \Lab_UT.S_0_s_axb3_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.S_0_s_axb3_LC_7_15_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.S_0_s_axb3_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(N__5633),
            .in2(_gnd_net_),
            .in3(N__5721),
            .lcout(\Lab_UT.S_0_s_axbZ0Z3 ),
            .ltout(\Lab_UT.S_0_s_axbZ0Z3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.S_m_am_3_LC_7_15_1 .C_ON=1'b0;
    defparam \Lab_UT.S_m_am_3_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.S_m_am_3_LC_7_15_1 .LUT_INIT=16'b0001111001111000;
    LogicCell40 \Lab_UT.S_m_am_3_LC_7_15_1  (
            .in0(N__5784),
            .in1(N__5863),
            .in2(N__3058),
            .in3(N__4635),
            .lcout(\Lab_UT.S_m_amZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.g1_2_LC_7_15_2 .C_ON=1'b0;
    defparam \Lab_UT.g1_2_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.g1_2_LC_7_15_2 .LUT_INIT=16'b1000101001000101;
    LogicCell40 \Lab_UT.g1_2_LC_7_15_2  (
            .in0(N__4397),
            .in1(N__4596),
            .in2(N__4489),
            .in3(N__4547),
            .lcout(\Lab_UT.g1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.gl_fsm.state_RNITO9T5_0_LC_7_15_3 .C_ON=1'b0;
    defparam \Glue_Lab2.gl_fsm.state_RNITO9T5_0_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.gl_fsm.state_RNITO9T5_0_LC_7_15_3 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \Glue_Lab2.gl_fsm.state_RNITO9T5_0_LC_7_15_3  (
            .in0(N__3535),
            .in1(N__4699),
            .in2(N__6361),
            .in3(N__5031),
            .lcout(\Glue_Lab2.Gl_r27_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.g0_4_1_LC_7_15_4 .C_ON=1'b0;
    defparam \Lab_UT.g0_4_1_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.g0_4_1_LC_7_15_4 .LUT_INIT=16'b0001001001001000;
    LogicCell40 \Lab_UT.g0_4_1_LC_7_15_4  (
            .in0(N__5864),
            .in1(N__5632),
            .in2(N__5811),
            .in3(N__5722),
            .lcout(\Lab_UT.g0_4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.S_m_bm_N_6L10_LC_7_15_5 .C_ON=1'b0;
    defparam \Lab_UT.S_m_bm_N_6L10_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.S_m_bm_N_6L10_LC_7_15_5 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \Lab_UT.S_m_bm_N_6L10_LC_7_15_5  (
            .in0(N__3559),
            .in1(N__4528),
            .in2(N__3580),
            .in3(N__4396),
            .lcout(\Lab_UT.S_m_bm_N_6LZ0Z10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.gl_fsm.state_RNITO9T5_0_0_LC_7_15_6 .C_ON=1'b0;
    defparam \Glue_Lab2.gl_fsm.state_RNITO9T5_0_0_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.gl_fsm.state_RNITO9T5_0_0_LC_7_15_6 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \Glue_Lab2.gl_fsm.state_RNITO9T5_0_0_LC_7_15_6  (
            .in0(N__4698),
            .in1(N__6348),
            .in2(N__5037),
            .in3(N__3534),
            .lcout(\Glue_Lab2.Gl_r17_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.S_0_s_c2_LC_7_15_7 .C_ON=1'b0;
    defparam \Lab_UT.S_0_s_c2_LC_7_15_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.S_0_s_c2_LC_7_15_7 .LUT_INIT=16'b1110110010000000;
    LogicCell40 \Lab_UT.S_0_s_c2_LC_7_15_7  (
            .in0(N__3558),
            .in1(N__4527),
            .in2(N__3579),
            .in3(N__4395),
            .lcout(\Lab_UT.S_0_s_cZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_r2_fast_0_LC_7_16_0 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_r2_fast_0_LC_7_16_0 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.Gl_r2_fast_0_LC_7_16_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Glue_Lab2.Gl_r2_fast_0_LC_7_16_0  (
            .in0(_gnd_net_),
            .in1(N__5388),
            .in2(_gnd_net_),
            .in3(N__6358),
            .lcout(Glue_Lab2_Gl_r2_fast_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6188),
            .ce(N__3627),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_r2_fast_2_LC_7_16_1 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_r2_fast_2_LC_7_16_1 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.Gl_r2_fast_2_LC_7_16_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Glue_Lab2.Gl_r2_fast_2_LC_7_16_1  (
            .in0(_gnd_net_),
            .in1(N__5227),
            .in2(_gnd_net_),
            .in3(N__6357),
            .lcout(Gl_r2_fast_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6188),
            .ce(N__3627),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_r2_2_rep1_LC_7_16_2 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_r2_2_rep1_LC_7_16_2 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.Gl_r2_2_rep1_LC_7_16_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Glue_Lab2.Gl_r2_2_rep1_LC_7_16_2  (
            .in0(N__6355),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5228),
            .lcout(Gl_r2_2_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6188),
            .ce(N__3627),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_r2_3_LC_7_16_3 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_r2_3_LC_7_16_3 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.Gl_r2_3_LC_7_16_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Glue_Lab2.Gl_r2_3_LC_7_16_3  (
            .in0(_gnd_net_),
            .in1(N__6356),
            .in2(_gnd_net_),
            .in3(N__6619),
            .lcout(Gl_r2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6188),
            .ce(N__3627),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_r2_0_LC_7_16_5 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_r2_0_LC_7_16_5 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.Gl_r2_0_LC_7_16_5 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \Glue_Lab2.Gl_r2_0_LC_7_16_5  (
            .in0(N__5389),
            .in1(N__6354),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(Gl_r2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6188),
            .ce(N__3627),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.de0.g0_LC_8_9_0 .C_ON=1'b0;
    defparam \Glue_Lab2.de0.g0_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.de0.g0_LC_8_9_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Glue_Lab2.de0.g0_LC_8_9_0  (
            .in0(N__5229),
            .in1(N__5439),
            .in2(N__3229),
            .in3(N__5387),
            .lcout(),
            .ltout(\Glue_Lab2.g0_9_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.reset_count_RNO_0_2_LC_8_9_1 .C_ON=1'b0;
    defparam \Glue_Lab2.reset_count_RNO_0_2_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.reset_count_RNO_0_2_LC_8_9_1 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \Glue_Lab2.reset_count_RNO_0_2_LC_8_9_1  (
            .in0(N__4198),
            .in1(N__5305),
            .in2(N__3151),
            .in3(N__3142),
            .lcout(\Glue_Lab2.reset_counte_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.de0.g0_4_LC_8_9_3 .C_ON=1'b0;
    defparam \Glue_Lab2.de0.g0_4_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.de0.g0_4_LC_8_9_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Glue_Lab2.de0.g0_4_LC_8_9_3  (
            .in0(N__4117),
            .in1(N__3848),
            .in2(N__4181),
            .in3(N__4032),
            .lcout(\Glue_Lab2.g0_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.de0.g0_0_LC_8_9_5 .C_ON=1'b0;
    defparam \Glue_Lab2.de0.g0_0_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.de0.g0_0_LC_8_9_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Glue_Lab2.de0.g0_0_LC_8_9_5  (
            .in0(N__4119),
            .in1(N__3849),
            .in2(N__4182),
            .in3(N__4034),
            .lcout(\Glue_Lab2.g0_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.de0.g0_12_LC_8_9_6 .C_ON=1'b0;
    defparam \Glue_Lab2.de0.g0_12_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.de0.g0_12_LC_8_9_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Glue_Lab2.de0.g0_12_LC_8_9_6  (
            .in0(N__4033),
            .in1(N__4118),
            .in2(N__4183),
            .in3(N__3852),
            .lcout(\Glue_Lab2.g0_7_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_4_LC_8_10_1 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_4_LC_8_10_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.bitcount_4_LC_8_10_1 .LUT_INIT=16'b1110111100100000;
    LogicCell40 \buart.Z_rx.bitcount_4_LC_8_10_1  (
            .in0(N__4178),
            .in1(N__3907),
            .in2(N__3970),
            .in3(N__3760),
            .lcout(buart__rx_bitcount_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6169),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNILM873_0_LC_8_10_2 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNILM873_0_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNILM873_0_LC_8_10_2 .LUT_INIT=16'b0000000011011111;
    LogicCell40 \buart.Z_rx.bitcount_RNILM873_0_LC_8_10_2  (
            .in0(N__3317),
            .in1(N__4075),
            .in2(N__3292),
            .in3(N__4314),
            .lcout(\buart.Z_rx.bitcountlde_0 ),
            .ltout(\buart.Z_rx.bitcountlde_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_0_LC_8_10_3 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_0_LC_8_10_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.bitcount_0_LC_8_10_3 .LUT_INIT=16'b1110111100100000;
    LogicCell40 \buart.Z_rx.bitcount_0_LC_8_10_3  (
            .in0(N__5447),
            .in1(N__3906),
            .in2(N__3136),
            .in3(N__3091),
            .lcout(buart__rx_bitcount_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6169),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNIIU223_0_LC_8_10_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNIIU223_0_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNIIU223_0_LC_8_10_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \buart.Z_rx.bitcount_RNIIU223_0_LC_8_10_4  (
            .in0(_gnd_net_),
            .in1(N__4313),
            .in2(_gnd_net_),
            .in3(N__4074),
            .lcout(\buart.Z_rx.N_29_0_i ),
            .ltout(\buart.Z_rx.N_29_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNO_0_0_LC_8_10_5 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNO_0_0_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNO_0_0_LC_8_10_5 .LUT_INIT=16'b0000011011110110;
    LogicCell40 \buart.Z_rx.bitcount_RNO_0_0_LC_8_10_5  (
            .in0(N__3119),
            .in1(N__5443),
            .in2(N__3094),
            .in3(N__3905),
            .lcout(\buart.Z_rx.bitcount_lm_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.de0.g0_2_LC_8_10_6 .C_ON=1'b0;
    defparam \Glue_Lab2.de0.g0_2_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.de0.g0_2_LC_8_10_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Glue_Lab2.de0.g0_2_LC_8_10_6  (
            .in0(N__5099),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6091),
            .lcout(\Glue_Lab2.de0.g0_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_8_10_7 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_8_10_7 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_8_10_7 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_1_LC_8_10_7  (
            .in0(N__3193),
            .in1(N__3220),
            .in2(_gnd_net_),
            .in3(N__3908),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6169),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNIMK771_1_4_LC_8_11_0 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNIMK771_1_4_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNIMK771_1_4_LC_8_11_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \buart.Z_rx.bitcount_RNIMK771_1_4_LC_8_11_0  (
            .in0(N__4028),
            .in1(N__4115),
            .in2(N__4179),
            .in3(N__3844),
            .lcout(\buart.Z_rx.un1_sample_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.de0.g0_7_LC_8_11_1 .C_ON=1'b0;
    defparam \Glue_Lab2.de0.g0_7_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.de0.g0_7_LC_8_11_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Glue_Lab2.de0.g0_7_LC_8_11_1  (
            .in0(N__4116),
            .in1(N__4164),
            .in2(N__3856),
            .in3(N__4029),
            .lcout(\Glue_Lab2.g0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.de0.g0_14_LC_8_11_2 .C_ON=1'b0;
    defparam \Glue_Lab2.de0.g0_14_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.de0.g0_14_LC_8_11_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Glue_Lab2.de0.g0_14_LC_8_11_2  (
            .in0(_gnd_net_),
            .in1(N__5104),
            .in2(_gnd_net_),
            .in3(N__5499),
            .lcout(),
            .ltout(\Glue_Lab2.de0.g0_5_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.de0.g0_11_LC_8_11_3 .C_ON=1'b0;
    defparam \Glue_Lab2.de0.g0_11_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.de0.g0_11_LC_8_11_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Glue_Lab2.de0.g0_11_LC_8_11_3  (
            .in0(N__5436),
            .in1(N__5230),
            .in2(N__3175),
            .in3(N__5355),
            .lcout(),
            .ltout(\Glue_Lab2.g0_9_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.reset_count_RNO_0_0_LC_8_11_4 .C_ON=1'b0;
    defparam \Glue_Lab2.reset_count_RNO_0_0_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.reset_count_RNO_0_0_LC_8_11_4 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \Glue_Lab2.reset_count_RNO_0_0_LC_8_11_4  (
            .in0(N__5294),
            .in1(N__3802),
            .in2(N__3172),
            .in3(N__3169),
            .lcout(\Glue_Lab2.reset_counte_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNIMK771_0_4_LC_8_11_5 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNIMK771_0_4_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNIMK771_0_4_LC_8_11_5 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \buart.Z_rx.bitcount_RNIMK771_0_4_LC_8_11_5  (
            .in0(N__4114),
            .in1(N__4027),
            .in2(N__3855),
            .in3(N__4160),
            .lcout(),
            .ltout(\buart.Z_rx.bitcount_RNIMK771_0Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNI9F1H1_0_LC_8_11_6 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNI9F1H1_0_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNI9F1H1_0_LC_8_11_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \buart.Z_rx.bitcount_RNI9F1H1_0_LC_8_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3154),
            .in3(N__5435),
            .lcout(bu_rx_data_rdy),
            .ltout(bu_rx_data_rdy_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.de0.de_esc_LC_8_11_7 .C_ON=1'b0;
    defparam \Glue_Lab2.de0.de_esc_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.de0.de_esc_LC_8_11_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Glue_Lab2.de0.de_esc_LC_8_11_7  (
            .in0(N__4900),
            .in1(N__4189),
            .in2(N__3451),
            .in3(N__5356),
            .lcout(\Glue_Lab2.i_rst_char_detected ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNI6KE3_5_LC_8_12_0 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI6KE3_5_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI6KE3_5_LC_8_12_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNI6KE3_5_LC_8_12_0  (
            .in0(N__3249),
            .in1(N__3407),
            .in2(N__3391),
            .in3(N__3376),
            .lcout(\buart.Z_rx.ser_clk_2_0 ),
            .ltout(\buart.Z_rx.ser_clk_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNIC77M1_0_LC_8_12_1 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNIC77M1_0_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNIC77M1_0_LC_8_12_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \buart.Z_rx.bitcount_RNIC77M1_0_LC_8_12_1  (
            .in0(N__3352),
            .in1(N__3319),
            .in2(N__3343),
            .in3(N__5453),
            .lcout(\buart.Z_rx.sample ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.de0.un2_de_hexplus_3_x0_LC_8_12_2 .C_ON=1'b0;
    defparam \Glue_Lab2.de0.un2_de_hexplus_3_x0_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.de0.un2_de_hexplus_3_x0_LC_8_12_2 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \Glue_Lab2.de0.un2_de_hexplus_3_x0_LC_8_12_2  (
            .in0(N__4231),
            .in1(N__5196),
            .in2(N__6471),
            .in3(N__5344),
            .lcout(),
            .ltout(\Glue_Lab2.de0.un2_de_hexplus_3_xZ0Z0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.de0.un2_de_hexplus_3_ns_LC_8_12_3 .C_ON=1'b0;
    defparam \Glue_Lab2.de0.un2_de_hexplus_3_ns_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.de0.un2_de_hexplus_3_ns_LC_8_12_3 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \Glue_Lab2.de0.un2_de_hexplus_3_ns_LC_8_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3340),
            .in3(N__6090),
            .lcout(),
            .ltout(\Glue_Lab2.de0.un2_de_hexplus_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.de0.de_hexplus_LC_8_12_4 .C_ON=1'b0;
    defparam \Glue_Lab2.de0.de_hexplus_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.de0.de_hexplus_LC_8_12_4 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \Glue_Lab2.de0.de_hexplus_LC_8_12_4  (
            .in0(N__3796),
            .in1(N__4237),
            .in2(N__3337),
            .in3(N__4312),
            .lcout(\Glue_Lab2.is_hexplus ),
            .ltout(\Glue_Lab2.is_hexplus_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_tx_data_4_LC_8_12_5 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_tx_data_4_LC_8_12_5 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.Gl_tx_data_4_LC_8_12_5 .LUT_INIT=16'b1010111110101111;
    LogicCell40 \Glue_Lab2.Gl_tx_data_4_LC_8_12_5  (
            .in0(N__5500),
            .in1(_gnd_net_),
            .in2(N__3334),
            .in3(_gnd_net_),
            .lcout(Gl_tx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6174),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_8_12_6 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_8_12_6 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_8_12_6 .LUT_INIT=16'b0000000001010010;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_2_LC_8_12_6  (
            .in0(N__3320),
            .in1(N__3284),
            .in2(N__3258),
            .in3(N__3942),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6174),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.gl_fsm.state_RNIDFRT_0_LC_8_12_7 .C_ON=1'b0;
    defparam \Glue_Lab2.gl_fsm.state_RNIDFRT_0_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.gl_fsm.state_RNIDFRT_0_LC_8_12_7 .LUT_INIT=16'b0000001000100000;
    LogicCell40 \Glue_Lab2.gl_fsm.state_RNIDFRT_0_LC_8_12_7  (
            .in0(N__5345),
            .in1(N__3527),
            .in2(N__6469),
            .in3(N__5197),
            .lcout(\Glue_Lab2.gl_fsm.enOp_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.gl_fsm.state_1_LC_8_13_0 .C_ON=1'b0;
    defparam \Glue_Lab2.gl_fsm.state_1_LC_8_13_0 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.gl_fsm.state_1_LC_8_13_0 .LUT_INIT=16'b0000001100100000;
    LogicCell40 \Glue_Lab2.gl_fsm.state_1_LC_8_13_0  (
            .in0(N__5010),
            .in1(N__6249),
            .in2(N__3533),
            .in3(N__4696),
            .lcout(Glue_Lab2_gl_fsm_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6179),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.gl_fsm.state_ns_1_0__m1_LC_8_13_1 .C_ON=1'b0;
    defparam \Glue_Lab2.gl_fsm.state_ns_1_0__m1_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.gl_fsm.state_ns_1_0__m1_LC_8_13_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Glue_Lab2.gl_fsm.state_ns_1_0__m1_LC_8_13_1  (
            .in0(_gnd_net_),
            .in1(N__3522),
            .in2(_gnd_net_),
            .in3(N__5008),
            .lcout(),
            .ltout(\Glue_Lab2.gl_fsm.N_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.gl_fsm.state_0_LC_8_13_2 .C_ON=1'b0;
    defparam \Glue_Lab2.gl_fsm.state_0_LC_8_13_2 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.gl_fsm.state_0_LC_8_13_2 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \Glue_Lab2.gl_fsm.state_0_LC_8_13_2  (
            .in0(N__6248),
            .in1(N__4695),
            .in2(N__3538),
            .in3(N__4268),
            .lcout(Glue_Lab2_gl_fsm_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6179),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.g0_LC_8_13_3 .C_ON=1'b0;
    defparam \Lab_UT.g0_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.g0_LC_8_13_3 .LUT_INIT=16'b0100110011101100;
    LogicCell40 \Lab_UT.g0_LC_8_13_3  (
            .in0(N__5950),
            .in1(N__3586),
            .in2(N__4288),
            .in3(N__3496),
            .lcout(),
            .ltout(led_c_0_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_tx_data_6_LC_8_13_4 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_tx_data_6_LC_8_13_4 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.Gl_tx_data_6_LC_8_13_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \Glue_Lab2.Gl_tx_data_6_LC_8_13_4  (
            .in0(N__5009),
            .in1(_gnd_net_),
            .in2(N__3490),
            .in3(N__5130),
            .lcout(Gl_tx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6179),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.S_m_bm_N_2L1_LC_8_13_6 .C_ON=1'b0;
    defparam \Lab_UT.S_m_bm_N_2L1_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.S_m_bm_N_2L1_LC_8_13_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.S_m_bm_N_2L1_LC_8_13_6  (
            .in0(_gnd_net_),
            .in1(N__5800),
            .in2(_gnd_net_),
            .in3(N__5873),
            .lcout(\Lab_UT.S_m_bm_N_2LZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.S_m_0_LC_8_13_7 .C_ON=1'b0;
    defparam \Lab_UT.S_m_0_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.S_m_0_LC_8_13_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \Lab_UT.S_m_0_LC_8_13_7  (
            .in0(N__4601),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4485),
            .lcout(led_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.S_1_ac0_1_0_0_LC_8_14_0 .C_ON=1'b0;
    defparam \Lab_UT.S_1_ac0_1_0_0_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.S_1_ac0_1_0_0_LC_8_14_0 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \Lab_UT.S_1_ac0_1_0_0_LC_8_14_0  (
            .in0(N__5805),
            .in1(N__4401),
            .in2(N__4558),
            .in3(N__5872),
            .lcout(\Lab_UT.S_1_ac0_1_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.S_1_axb1_LC_8_14_1 .C_ON=1'b0;
    defparam \Lab_UT.S_1_axb1_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.S_1_axb1_LC_8_14_1 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \Lab_UT.S_1_axb1_LC_8_14_1  (
            .in0(N__4402),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4556),
            .lcout(),
            .ltout(\Lab_UT.S_1_axbZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.S_1_ac0_1_0_LC_8_14_2 .C_ON=1'b0;
    defparam \Lab_UT.S_1_ac0_1_0_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.S_1_ac0_1_0_LC_8_14_2 .LUT_INIT=16'b1110110011111100;
    LogicCell40 \Lab_UT.S_1_ac0_1_0_LC_8_14_2  (
            .in0(N__4595),
            .in1(N__3610),
            .in2(N__3604),
            .in3(N__4478),
            .lcout(\Lab_UT.S_1_c3_d ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.S_m_am_1_LC_8_14_3 .C_ON=1'b0;
    defparam \Lab_UT.S_m_am_1_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.S_m_am_1_LC_8_14_3 .LUT_INIT=16'b1001010101101010;
    LogicCell40 \Lab_UT.S_m_am_1_LC_8_14_3  (
            .in0(N__4400),
            .in1(N__4594),
            .in2(N__4487),
            .in3(N__4552),
            .lcout(\Lab_UT.S_m_amZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_r1_0_LC_8_14_4 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_r1_0_LC_8_14_4 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.Gl_r1_0_LC_8_14_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Glue_Lab2.Gl_r1_0_LC_8_14_4  (
            .in0(_gnd_net_),
            .in1(N__6291),
            .in2(_gnd_net_),
            .in3(N__5383),
            .lcout(Gl_r1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6185),
            .ce(N__3673),
            .sr(_gnd_net_));
    defparam \Lab_UT.g1_0_LC_8_14_5 .C_ON=1'b0;
    defparam \Lab_UT.g1_0_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.g1_0_LC_8_14_5 .LUT_INIT=16'b1000101001000101;
    LogicCell40 \Lab_UT.g1_0_LC_8_14_5  (
            .in0(N__4398),
            .in1(N__4590),
            .in2(N__4486),
            .in3(N__4550),
            .lcout(\Lab_UT.g1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.g0_7_LC_8_14_6 .C_ON=1'b0;
    defparam \Lab_UT.g0_7_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.g0_7_LC_8_14_6 .LUT_INIT=16'b1110100010001000;
    LogicCell40 \Lab_UT.g0_7_LC_8_14_6  (
            .in0(N__4551),
            .in1(N__4399),
            .in2(N__4602),
            .in3(N__4474),
            .lcout(),
            .ltout(\Lab_UT.S_0_s_c2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.g1_LC_8_14_7 .C_ON=1'b0;
    defparam \Lab_UT.g1_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.g1_LC_8_14_7 .LUT_INIT=16'b1111111111000000;
    LogicCell40 \Lab_UT.g1_LC_8_14_7  (
            .in0(_gnd_net_),
            .in1(N__3679),
            .in2(N__3595),
            .in3(N__3592),
            .lcout(\Lab_UT.gZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.S_m_bm_1_2_LC_8_15_0 .C_ON=1'b0;
    defparam \Lab_UT.S_m_bm_1_2_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.S_m_bm_1_2_LC_8_15_0 .LUT_INIT=16'b0100110101000100;
    LogicCell40 \Lab_UT.S_m_bm_1_2_LC_8_15_0  (
            .in0(N__4394),
            .in1(N__4526),
            .in2(N__3557),
            .in3(N__3572),
            .lcout(\Lab_UT.S_m_bm_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_r1_fast_0_LC_8_15_1 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_r1_fast_0_LC_8_15_1 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.Gl_r1_fast_0_LC_8_15_1 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \Glue_Lab2.Gl_r1_fast_0_LC_8_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6359),
            .in3(N__5386),
            .lcout(Glue_Lab2_Gl_r1_fast_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6189),
            .ce(N__3672),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_r1_fast_2_LC_8_15_2 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_r1_fast_2_LC_8_15_2 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.Gl_r1_fast_2_LC_8_15_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \Glue_Lab2.Gl_r1_fast_2_LC_8_15_2  (
            .in0(N__5234),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6343),
            .lcout(Gl_r1_fast_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6189),
            .ce(N__3672),
            .sr(_gnd_net_));
    defparam \Lab_UT.S_m_bm_N_5L7_LC_8_15_3 .C_ON=1'b0;
    defparam \Lab_UT.S_m_bm_N_5L7_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.S_m_bm_N_5L7_LC_8_15_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \Lab_UT.S_m_bm_N_5L7_LC_8_15_3  (
            .in0(N__4746),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4734),
            .lcout(\Lab_UT.S_m_bm_N_5LZ0Z7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_r1_2_rep1_LC_8_15_4 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_r1_2_rep1_LC_8_15_4 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.Gl_r1_2_rep1_LC_8_15_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \Glue_Lab2.Gl_r1_2_rep1_LC_8_15_4  (
            .in0(N__5233),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6339),
            .lcout(Gl_r1_2_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6189),
            .ce(N__3672),
            .sr(_gnd_net_));
    defparam \Lab_UT.g0_4_0_LC_8_15_5 .C_ON=1'b0;
    defparam \Lab_UT.g0_4_0_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.g0_4_0_LC_8_15_5 .LUT_INIT=16'b0001001001001000;
    LogicCell40 \Lab_UT.g0_4_0_LC_8_15_5  (
            .in0(N__3727),
            .in1(N__5631),
            .in2(N__3705),
            .in3(N__5723),
            .lcout(\Lab_UT.g0_4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_r1_2_LC_8_15_6 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_r1_2_LC_8_15_6 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.Gl_r1_2_LC_8_15_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \Glue_Lab2.Gl_r1_2_LC_8_15_6  (
            .in0(N__5232),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6338),
            .lcout(Gl_r1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6189),
            .ce(N__3672),
            .sr(_gnd_net_));
    defparam \Lab_UT.g0_4_LC_8_15_7 .C_ON=1'b0;
    defparam \Lab_UT.g0_4_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.g0_4_LC_8_15_7 .LUT_INIT=16'b1110110010000000;
    LogicCell40 \Lab_UT.g0_4_LC_8_15_7  (
            .in0(N__5860),
            .in1(N__5630),
            .in2(N__5801),
            .in3(N__5724),
            .lcout(\Lab_UT.S_0_s_ac0_5_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.g0_1_1_LC_8_16_0 .C_ON=1'b0;
    defparam \Lab_UT.g0_1_1_LC_8_16_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.g0_1_1_LC_8_16_0 .LUT_INIT=16'b0011101100001010;
    LogicCell40 \Lab_UT.g0_1_1_LC_8_16_0  (
            .in0(N__5871),
            .in1(N__4546),
            .in2(N__5812),
            .in3(N__4416),
            .lcout(\Lab_UT.g0_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_r2_1_LC_8_16_1 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_r2_1_LC_8_16_1 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.Gl_r2_1_LC_8_16_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Glue_Lab2.Gl_r2_1_LC_8_16_1  (
            .in0(_gnd_net_),
            .in1(N__6344),
            .in2(_gnd_net_),
            .in3(N__6475),
            .lcout(Gl_r2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6192),
            .ce(N__3628),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_r2_2_LC_8_16_2 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_r2_2_LC_8_16_2 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.Gl_r2_2_LC_8_16_2 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \Glue_Lab2.Gl_r2_2_LC_8_16_2  (
            .in0(N__5235),
            .in1(_gnd_net_),
            .in2(N__6360),
            .in3(_gnd_net_),
            .lcout(Gl_r2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6192),
            .ce(N__3628),
            .sr(_gnd_net_));
    defparam \Lab_UT.g0_2_LC_8_16_3 .C_ON=1'b0;
    defparam \Lab_UT.g0_2_LC_8_16_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.g0_2_LC_8_16_3 .LUT_INIT=16'b1110100010100000;
    LogicCell40 \Lab_UT.g0_2_LC_8_16_3  (
            .in0(N__4415),
            .in1(N__4449),
            .in2(N__4557),
            .in3(N__4603),
            .lcout(),
            .ltout(\Lab_UT.S_0_s_c2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.g1_1_LC_8_16_4 .C_ON=1'b0;
    defparam \Lab_UT.g1_1_LC_8_16_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.g1_1_LC_8_16_4 .LUT_INIT=16'b1111111111000000;
    LogicCell40 \Lab_UT.g1_1_LC_8_16_4  (
            .in0(_gnd_net_),
            .in1(N__3616),
            .in2(N__3790),
            .in3(N__3787),
            .lcout(Lab_UT_g1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_9_9_0 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_9_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_c_0_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(N__5438),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(\buart.Z_rx.bitcount_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_9_9_1 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_9_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(N__4035),
            .in2(_gnd_net_),
            .in3(N__3772),
            .lcout(\buart.Z_rx.bitcount_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_0 ),
            .carryout(\buart.Z_rx.bitcount_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_9_9_2 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_9_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(N__3853),
            .in2(_gnd_net_),
            .in3(N__3769),
            .lcout(\buart.Z_rx.bitcount_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_1 ),
            .carryout(\buart.Z_rx.bitcount_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_9_9_3 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_9_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_9_9_3  (
            .in0(_gnd_net_),
            .in1(N__4122),
            .in2(_gnd_net_),
            .in3(N__3766),
            .lcout(\buart.Z_rx.bitcount_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_2 ),
            .carryout(\buart.Z_rx.bitcount_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNO_0_4_LC_9_9_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNO_0_4_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNO_0_4_LC_9_9_4 .LUT_INIT=16'b0001101101001110;
    LogicCell40 \buart.Z_rx.bitcount_RNO_0_4_LC_9_9_4  (
            .in0(N__3985),
            .in1(N__4177),
            .in2(N__3928),
            .in3(N__3763),
            .lcout(\buart.Z_rx.bitcount_lm_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNO_0_1_LC_9_9_7 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNO_0_1_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNO_0_1_LC_9_9_7 .LUT_INIT=16'b0000111101100110;
    LogicCell40 \buart.Z_rx.bitcount_RNO_0_1_LC_9_9_7  (
            .in0(N__3754),
            .in1(N__4036),
            .in2(N__3927),
            .in3(N__3986),
            .lcout(\buart.Z_rx.bitcount_lm_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNO_0_3_LC_9_10_0 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNO_0_3_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNO_0_3_LC_9_10_0 .LUT_INIT=16'b0000111101100110;
    LogicCell40 \buart.Z_rx.bitcount_RNO_0_3_LC_9_10_0  (
            .in0(N__4123),
            .in1(N__3748),
            .in2(N__3941),
            .in3(N__3988),
            .lcout(),
            .ltout(\buart.Z_rx.bitcount_lm_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_3_LC_9_10_1 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_3_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.bitcount_3_LC_9_10_1 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \buart.Z_rx.bitcount_3_LC_9_10_1  (
            .in0(N__4121),
            .in1(N__3969),
            .in2(N__3742),
            .in3(N__3923),
            .lcout(buart__rx_bitcount_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6171),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNIMK771_4_LC_9_10_2 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNIMK771_4_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNIMK771_4_LC_9_10_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \buart.Z_rx.bitcount_RNIMK771_4_LC_9_10_2  (
            .in0(N__3850),
            .in1(N__4030),
            .in2(N__4180),
            .in3(N__4120),
            .lcout(),
            .ltout(\buart.Z_rx.bitcount_RNIMK771Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNI9F1H1_0_0_LC_9_10_3 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNI9F1H1_0_0_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNI9F1H1_0_0_LC_9_10_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \buart.Z_rx.bitcount_RNI9F1H1_0_0_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4078),
            .in3(N__5437),
            .lcout(\buart.Z_rx.idle ),
            .ltout(\buart.Z_rx.idle_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.hh_RNI065O1_0_LC_9_10_4 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_RNI065O1_0_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.hh_RNI065O1_0_LC_9_10_4 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \buart.Z_rx.hh_RNI065O1_0_LC_9_10_4  (
            .in0(_gnd_net_),
            .in1(N__4218),
            .in2(N__4066),
            .in3(N__4063),
            .lcout(\buart.Z_rx.startbit ),
            .ltout(\buart.Z_rx.startbit_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_1_LC_9_10_5 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_1_LC_9_10_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.bitcount_1_LC_9_10_5 .LUT_INIT=16'b1111101100001000;
    LogicCell40 \buart.Z_rx.bitcount_1_LC_9_10_5  (
            .in0(N__4031),
            .in1(N__3967),
            .in2(N__4045),
            .in3(N__4042),
            .lcout(buart__rx_bitcount_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6171),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNO_0_2_LC_9_10_6 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNO_0_2_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNO_0_2_LC_9_10_6 .LUT_INIT=16'b0000111101100110;
    LogicCell40 \buart.Z_rx.bitcount_RNO_0_2_LC_9_10_6  (
            .in0(N__3851),
            .in1(N__3994),
            .in2(N__3940),
            .in3(N__3987),
            .lcout(),
            .ltout(\buart.Z_rx.bitcount_lm_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_2_LC_9_10_7 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_2_LC_9_10_7 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.bitcount_2_LC_9_10_7 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \buart.Z_rx.bitcount_2_LC_9_10_7  (
            .in0(N__3854),
            .in1(N__3968),
            .in2(N__3949),
            .in3(N__3922),
            .lcout(buart__rx_bitcount_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6171),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.de0.g0_13_LC_9_11_0 .C_ON=1'b0;
    defparam \Glue_Lab2.de0.g0_13_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.de0.g0_13_LC_9_11_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Glue_Lab2.de0.g0_13_LC_9_11_0  (
            .in0(N__6659),
            .in1(N__6446),
            .in2(N__6535),
            .in3(N__6576),
            .lcout(\Glue_Lab2.g0_8_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_3_LC_9_11_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_3_LC_9_11_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.shifter_3_LC_9_11_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_3_LC_9_11_1  (
            .in0(N__5495),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6175),
            .ce(N__6073),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.de0.un2_de_hexplus_2_LC_9_11_2 .C_ON=1'b0;
    defparam \Glue_Lab2.de0.un2_de_hexplus_2_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.de0.un2_de_hexplus_2_LC_9_11_2 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \Glue_Lab2.de0.un2_de_hexplus_2_LC_9_11_2  (
            .in0(N__5101),
            .in1(_gnd_net_),
            .in2(N__6673),
            .in3(N__6572),
            .lcout(\Glue_Lab2.de0.un2_de_hexplusZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_6_LC_9_11_3 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_6_LC_9_11_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.shifter_6_LC_9_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_6_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6660),
            .lcout(bu_rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6175),
            .ce(N__6073),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.de0.un1_charData_LC_9_11_4 .C_ON=1'b0;
    defparam \Glue_Lab2.de0.un1_charData_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.de0.un1_charData_LC_9_11_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Glue_Lab2.de0.un1_charData_LC_9_11_4  (
            .in0(N__5100),
            .in1(N__4230),
            .in2(N__6672),
            .in3(N__5493),
            .lcout(\Glue_Lab2.de0.un1_charDataZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_fast_5_LC_9_11_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_5_LC_9_11_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.shifter_fast_5_LC_9_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_fast_5_LC_9_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5103),
            .lcout(buart__rx_shifter_fast_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6175),
            .ce(N__6073),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_7_LC_9_11_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_7_LC_9_11_6 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.shifter_7_LC_9_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_7_LC_9_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4219),
            .lcout(bu_rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6175),
            .ce(N__6073),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.gl_fsm.enOp_0_a2_4_LC_9_11_7 .C_ON=1'b0;
    defparam \Glue_Lab2.gl_fsm.enOp_0_a2_4_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.gl_fsm.enOp_0_a2_4_LC_9_11_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Glue_Lab2.gl_fsm.enOp_0_a2_4_LC_9_11_7  (
            .in0(N__5494),
            .in1(N__6530),
            .in2(N__6595),
            .in3(N__5102),
            .lcout(\Glue_Lab2.gl_fsm.enOp_0_a2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.de0.g0_1_LC_9_12_0 .C_ON=1'b0;
    defparam \Glue_Lab2.de0.g0_1_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.de0.g0_1_LC_9_12_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Glue_Lab2.de0.g0_1_LC_9_12_0  (
            .in0(N__6662),
            .in1(N__6578),
            .in2(N__6534),
            .in3(N__6460),
            .lcout(\Glue_Lab2.g0_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_1_LC_9_12_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_1_LC_9_12_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.shifter_1_LC_9_12_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \buart.Z_rx.shifter_1_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(N__5226),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6180),
            .ce(N__6058),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.de0.de_esc_3_LC_9_12_2 .C_ON=1'b0;
    defparam \Glue_Lab2.de0.de_esc_3_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.de0.de_esc_3_LC_9_12_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Glue_Lab2.de0.de_esc_3_LC_9_12_2  (
            .in0(N__6661),
            .in1(N__6577),
            .in2(_gnd_net_),
            .in3(N__6461),
            .lcout(\Glue_Lab2.de0.de_escZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_0_LC_9_12_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_LC_9_12_6 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.shifter_0_LC_9_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_LC_9_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6462),
            .lcout(bu_rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6180),
            .ce(N__6058),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.gl_fsm.state_RNIQ3DV3_0_LC_9_12_7 .C_ON=1'b0;
    defparam \Glue_Lab2.gl_fsm.state_RNIQ3DV3_0_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.gl_fsm.state_RNIQ3DV3_0_LC_9_12_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Glue_Lab2.gl_fsm.state_RNIQ3DV3_0_LC_9_12_7  (
            .in0(N__4666),
            .in1(N__4330),
            .in2(N__4324),
            .in3(N__4315),
            .lcout(\Glue_Lab2.enOp ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_rst_RNI7BQG_LC_9_13_0 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_rst_RNI7BQG_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.Gl_rst_RNI7BQG_LC_9_13_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Glue_Lab2.Gl_rst_RNI7BQG_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(N__6450),
            .in2(_gnd_net_),
            .in3(N__6309),
            .lcout(),
            .ltout(\Glue_Lab2.Gl_r1_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_Op_1_LC_9_13_1 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_Op_1_LC_9_13_1 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.Gl_Op_1_LC_9_13_1 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \Glue_Lab2.Gl_Op_1_LC_9_13_1  (
            .in0(N__5977),
            .in1(N__6337),
            .in2(N__4294),
            .in3(N__4274),
            .lcout(Glue_Lab2_Gl_Op_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6186),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_rst_RNI8CQG_LC_9_13_2 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_rst_RNI8CQG_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.Gl_rst_RNI8CQG_LC_9_13_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Glue_Lab2.Gl_rst_RNI8CQG_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(N__6310),
            .in2(_gnd_net_),
            .in3(N__5231),
            .lcout(),
            .ltout(\Glue_Lab2.Gl_r1_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_Op_2_LC_9_13_3 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_Op_2_LC_9_13_3 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.Gl_Op_2_LC_9_13_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \Glue_Lab2.Gl_Op_2_LC_9_13_3  (
            .in0(N__6311),
            .in1(N__4275),
            .in2(N__4291),
            .in3(N__5916),
            .lcout(Glue_Lab2_Gl_Op_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6186),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_Op_5_LC_9_13_4 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_Op_5_LC_9_13_4 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.Gl_Op_5_LC_9_13_4 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \Glue_Lab2.Gl_Op_5_LC_9_13_4  (
            .in0(N__4273),
            .in1(N__6313),
            .in2(_gnd_net_),
            .in3(N__5951),
            .lcout(Glue_Lab2_Gl_Op_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6186),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.g0_1_2_LC_9_13_5 .C_ON=1'b0;
    defparam \Lab_UT.g0_1_2_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.g0_1_2_LC_9_13_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \Lab_UT.g0_1_2_LC_9_13_5  (
            .in0(N__6029),
            .in1(N__6005),
            .in2(N__5982),
            .in3(N__5915),
            .lcout(\Lab_UT.g0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_Op_3_LC_9_13_6 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_Op_3_LC_9_13_6 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.Gl_Op_3_LC_9_13_6 .LUT_INIT=16'b0000000011111010;
    LogicCell40 \Glue_Lab2.Gl_Op_3_LC_9_13_6  (
            .in0(N__6006),
            .in1(_gnd_net_),
            .in2(N__4276),
            .in3(N__6312),
            .lcout(Glue_Lab2_Gl_Op_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6186),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_Op_0_LC_9_13_7 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_Op_0_LC_9_13_7 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.Gl_Op_0_LC_9_13_7 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \Glue_Lab2.Gl_Op_0_LC_9_13_7  (
            .in0(N__6030),
            .in1(N__6336),
            .in2(_gnd_net_),
            .in3(N__4269),
            .lcout(Glue_Lab2_Gl_Op_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6186),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_tx_data_2_LC_9_14_0 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_tx_data_2_LC_9_14_0 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.Gl_tx_data_2_LC_9_14_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Glue_Lab2.Gl_tx_data_2_LC_9_14_0  (
            .in0(N__4614),
            .in1(N__5032),
            .in2(_gnd_net_),
            .in3(N__5236),
            .lcout(Gl_tx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6190),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.gl_fsm.state_RNIIM7B_1_LC_9_14_3 .C_ON=1'b0;
    defparam \Glue_Lab2.gl_fsm.state_RNIIM7B_1_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.gl_fsm.state_RNIIM7B_1_LC_9_14_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Glue_Lab2.gl_fsm.state_RNIIM7B_1_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(N__4689),
            .in2(_gnd_net_),
            .in3(N__6674),
            .lcout(\Glue_Lab2.gl_fsm.enOp_0_a2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_Op_RNIDA8P_2_LC_9_14_5 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_Op_RNIDA8P_2_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.Gl_Op_RNIDA8P_2_LC_9_14_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Glue_Lab2.Gl_Op_RNIDA8P_2_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(N__6001),
            .in2(_gnd_net_),
            .in3(N__5914),
            .lcout(),
            .ltout(\Glue_Lab2.Gl_subtract_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_Op_RNIFO4V1_0_LC_9_14_6 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_Op_RNIFO4V1_0_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.Gl_Op_RNIFO4V1_0_LC_9_14_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Glue_Lab2.Gl_Op_RNIFO4V1_0_LC_9_14_6  (
            .in0(N__5952),
            .in1(N__5981),
            .in2(N__4657),
            .in3(N__6025),
            .lcout(Gl_subtract),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.S_0_s_ac0_5_d_LC_9_15_0 .C_ON=1'b0;
    defparam \Lab_UT.S_0_s_ac0_5_d_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.S_0_s_ac0_5_d_LC_9_15_0 .LUT_INIT=16'b0100000010000000;
    LogicCell40 \Lab_UT.S_0_s_ac0_5_d_LC_9_15_0  (
            .in0(N__5862),
            .in1(N__4654),
            .in2(N__4645),
            .in3(N__5780),
            .lcout(\Lab_UT.S_0_s_ac0_5_dZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.S_m_am_2_LC_9_15_3 .C_ON=1'b0;
    defparam \Lab_UT.S_m_am_2_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.S_m_am_2_LC_9_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Lab_UT.S_m_am_2_LC_9_15_3  (
            .in0(N__5779),
            .in1(N__5861),
            .in2(_gnd_net_),
            .in3(N__4641),
            .lcout(),
            .ltout(\Lab_UT.S_m_amZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.S_m_ns_2_LC_9_15_4 .C_ON=1'b0;
    defparam \Lab_UT.S_m_ns_2_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.S_m_ns_2_LC_9_15_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \Lab_UT.S_m_ns_2_LC_9_15_4  (
            .in0(_gnd_net_),
            .in1(N__4717),
            .in2(N__4624),
            .in3(N__5557),
            .lcout(led_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.S_m_bm_1_LC_9_15_5 .C_ON=1'b0;
    defparam \Lab_UT.S_m_bm_1_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.S_m_bm_1_LC_9_15_5 .LUT_INIT=16'b0110001110011100;
    LogicCell40 \Lab_UT.S_m_bm_1_LC_9_15_5  (
            .in0(N__4597),
            .in1(N__4548),
            .in2(N__4488),
            .in3(N__4420),
            .lcout(),
            .ltout(\Lab_UT.S_m_bmZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.S_m_ns_1_LC_9_15_6 .C_ON=1'b0;
    defparam \Lab_UT.S_m_ns_1_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.S_m_ns_1_LC_9_15_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \Lab_UT.S_m_ns_1_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(N__4351),
            .in2(N__4345),
            .in3(N__5558),
            .lcout(led_c_1),
            .ltout(led_c_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_tx_data_1_LC_9_15_7 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_tx_data_1_LC_9_15_7 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.Gl_tx_data_1_LC_9_15_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \Glue_Lab2.Gl_tx_data_1_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(N__6470),
            .in2(N__4765),
            .in3(N__5033),
            .lcout(Gl_tx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6193),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.S_m_bm_2_LC_9_16_1 .C_ON=1'b0;
    defparam \Lab_UT.S_m_bm_2_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.S_m_bm_2_LC_9_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Lab_UT.S_m_bm_2_LC_9_16_1  (
            .in0(N__4750),
            .in1(N__4735),
            .in2(_gnd_net_),
            .in3(N__4723),
            .lcout(\Lab_UT.S_m_bmZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNI1O14_1_LC_11_7_0 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI1O14_1_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI1O14_1_LC_11_7_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNI1O14_1_LC_11_7_0  (
            .in0(_gnd_net_),
            .in1(N__4839),
            .in2(_gnd_net_),
            .in3(N__4817),
            .lcout(\buart.Z_tx.Z_baudgen.un2_counter_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_11_7_1 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_11_7_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_11_7_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_0_LC_11_7_1  (
            .in0(N__4818),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6182),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_11_7_7 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_11_7_7 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_11_7_7 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_1_LC_11_7_7  (
            .in0(N__4819),
            .in1(_gnd_net_),
            .in2(N__4843),
            .in3(_gnd_net_),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6182),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_11_8_0 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_11_8_0 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_11_8_0 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_4_LC_11_8_0  (
            .in0(N__4888),
            .in1(N__6820),
            .in2(N__6886),
            .in3(N__6908),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6177),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNIQJ4A_4_LC_11_8_1 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIQJ4A_4_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIQJ4A_4_LC_11_8_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNIQJ4A_4_LC_11_8_1  (
            .in0(N__6907),
            .in1(N__4887),
            .in2(N__6823),
            .in3(N__6881),
            .lcout(\buart.Z_tx.Z_baudgen.un2_counter_c5 ),
            .ltout(\buart.Z_tx.Z_baudgen.un2_counter_c5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_11_8_2 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_11_8_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_11_8_2 .LUT_INIT=16'b0000000001011010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_5_LC_11_8_2  (
            .in0(N__4871),
            .in1(_gnd_net_),
            .in2(N__4711),
            .in3(N__6855),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6177),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNINP26_6_LC_11_8_3 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNINP26_6_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNINP26_6_LC_11_8_3 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNINP26_6_LC_11_8_3  (
            .in0(N__4853),
            .in1(N__4837),
            .in2(_gnd_net_),
            .in3(N__4815),
            .lcout(\buart.Z_tx.Z_baudgen.un1_bitcount_c2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_11_8_4 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_11_8_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_11_8_4 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_6_LC_11_8_4  (
            .in0(N__4872),
            .in1(N__4855),
            .in2(N__4708),
            .in3(N__6856),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6177),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNIES38_0_4_LC_11_8_5 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIES38_0_4_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIES38_0_4_LC_11_8_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNIES38_0_4_LC_11_8_5  (
            .in0(N__6906),
            .in1(N__4886),
            .in2(N__6822),
            .in3(N__4870),
            .lcout(\buart.Z_tx.Z_baudgen.counter_RNIES38_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNIES38_4_LC_11_8_6 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIES38_4_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIES38_4_LC_11_8_6 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNIES38_4_LC_11_8_6  (
            .in0(N__4885),
            .in1(N__6813),
            .in2(N__4873),
            .in3(N__6905),
            .lcout(),
            .ltout(\buart.Z_tx.Z_baudgen.ser_clk_sx_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_6_LC_11_8_7 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_6_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_6_LC_11_8_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNI5M6E_6_LC_11_8_7  (
            .in0(N__4854),
            .in1(N__4838),
            .in2(N__4822),
            .in3(N__4816),
            .lcout(\buart.Z_tx.ser_clk ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNIBADL_1_LC_11_9_0 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIBADL_1_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIBADL_1_LC_11_9_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \buart.Z_tx.bitcount_RNIBADL_1_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__4959),
            .in2(_gnd_net_),
            .in3(N__4919),
            .lcout(),
            .ltout(\buart.Z_tx.bitcount_RNIBADLZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNIVE1P1_4_LC_11_9_1 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIVE1P1_4_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIVE1P1_4_LC_11_9_1 .LUT_INIT=16'b0000001000100010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNIVE1P1_4_LC_11_9_1  (
            .in0(N__4798),
            .in1(N__4792),
            .in2(N__4786),
            .in3(N__4774),
            .lcout(\buart.Z_tx.counter_RNIVE1P1_4 ),
            .ltout(\buart.Z_tx.counter_RNIVE1P1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_2_LC_11_9_2 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_2_LC_11_9_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.bitcount_2_LC_11_9_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \buart.Z_tx.bitcount_2_LC_11_9_2  (
            .in0(N__6786),
            .in1(N__5068),
            .in2(N__4783),
            .in3(N__4780),
            .lcout(\buart.Z_tx.bitcountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6172),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_11_9_3 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_11_9_3 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \buart.Z_tx.bitcount_RNO_0_2_LC_11_9_3  (
            .in0(N__4921),
            .in1(N__4961),
            .in2(_gnd_net_),
            .in3(N__6848),
            .lcout(\buart.Z_tx.un1_bitcount_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNIFEDL_3_LC_11_9_4 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIFEDL_3_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIFEDL_3_LC_11_9_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \buart.Z_tx.bitcount_RNIFEDL_3_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(N__5052),
            .in2(_gnd_net_),
            .in3(N__5066),
            .lcout(\buart.Z_tx.uart_busy_0_0 ),
            .ltout(\buart.Z_tx.uart_busy_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNIQL5G1_1_LC_11_9_5 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIQL5G1_1_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIQL5G1_1_LC_11_9_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \buart.Z_tx.bitcount_RNIQL5G1_1_LC_11_9_5  (
            .in0(N__4920),
            .in1(N__6785),
            .in2(N__4768),
            .in3(N__4960),
            .lcout(\buart.Z_tx.un1_uart_wr_i_0_i_sx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_11_9_6 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_11_9_6 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \buart.Z_tx.bitcount_RNO_0_3_LC_11_9_6  (
            .in0(N__6849),
            .in1(N__4922),
            .in2(N__4966),
            .in3(N__5067),
            .lcout(),
            .ltout(\buart.Z_tx.un1_bitcount_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_3_LC_11_9_7 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_3_LC_11_9_7 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.bitcount_3_LC_11_9_7 .LUT_INIT=16'b1110110111011110;
    LogicCell40 \buart.Z_tx.bitcount_3_LC_11_9_7  (
            .in0(N__5053),
            .in1(N__6787),
            .in2(N__5056),
            .in3(N__4939),
            .lcout(\buart.Z_tx.bitcountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6172),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNIV8N32_1_LC_11_10_2 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIV8N32_1_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIV8N32_1_LC_11_10_2 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \buart.Z_tx.bitcount_RNIV8N32_1_LC_11_10_2  (
            .in0(N__6859),
            .in1(N__6761),
            .in2(_gnd_net_),
            .in3(N__5044),
            .lcout(\buart.Z_tx.un1_uart_wr_i_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_tx_data_rdy_LC_11_10_4 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_tx_data_rdy_LC_11_10_4 .SEQ_MODE=4'b1000;
    defparam \Glue_Lab2.Gl_tx_data_rdy_LC_11_10_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \Glue_Lab2.Gl_tx_data_rdy_LC_11_10_4  (
            .in0(N__6202),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5038),
            .lcout(Gl_tx_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6176),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNO_0_1_LC_11_10_5 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNO_0_1_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNO_0_1_LC_11_10_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \buart.Z_tx.bitcount_RNO_0_1_LC_11_10_5  (
            .in0(_gnd_net_),
            .in1(N__4923),
            .in2(_gnd_net_),
            .in3(N__6858),
            .lcout(),
            .ltout(\buart.Z_tx.un1_bitcount_c1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_1_LC_11_10_6 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_1_LC_11_10_6 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.bitcount_1_LC_11_10_6 .LUT_INIT=16'b1110110111011110;
    LogicCell40 \buart.Z_tx.bitcount_1_LC_11_10_6  (
            .in0(N__4938),
            .in1(N__6763),
            .in2(N__4969),
            .in3(N__4965),
            .lcout(\buart.Z_tx.bitcountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6176),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_0_LC_11_10_7 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_0_LC_11_10_7 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.bitcount_0_LC_11_10_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_tx.bitcount_0_LC_11_10_7  (
            .in0(N__6762),
            .in1(N__4924),
            .in2(_gnd_net_),
            .in3(N__4937),
            .lcout(\buart.Z_tx.bitcountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6176),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.de0.de_esc_4_LC_11_11_0 .C_ON=1'b0;
    defparam \Glue_Lab2.de0.de_esc_4_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.de0.de_esc_4_LC_11_11_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \Glue_Lab2.de0.de_esc_4_LC_11_11_0  (
            .in0(N__5487),
            .in1(N__6505),
            .in2(N__5129),
            .in3(N__5175),
            .lcout(\Glue_Lab2.de0.de_escZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.de0.g0_10_LC_11_11_1 .C_ON=1'b0;
    defparam \Glue_Lab2.de0.g0_10_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.de0.g0_10_LC_11_11_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Glue_Lab2.de0.g0_10_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(N__5118),
            .in2(_gnd_net_),
            .in3(N__5489),
            .lcout(),
            .ltout(\Glue_Lab2.de0.g0_5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.de0.g0_3_LC_11_11_2 .C_ON=1'b0;
    defparam \Glue_Lab2.de0.g0_3_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.de0.g0_3_LC_11_11_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Glue_Lab2.de0.g0_3_LC_11_11_2  (
            .in0(N__5454),
            .in1(N__5177),
            .in2(N__5527),
            .in3(N__5385),
            .lcout(),
            .ltout(\Glue_Lab2.g0_9_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.reset_count_RNO_0_1_LC_11_11_3 .C_ON=1'b0;
    defparam \Glue_Lab2.reset_count_RNO_0_1_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.reset_count_RNO_0_1_LC_11_11_3 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \Glue_Lab2.reset_count_RNO_0_1_LC_11_11_3  (
            .in0(N__5303),
            .in1(N__6388),
            .in2(N__5524),
            .in3(N__5521),
            .lcout(\Glue_Lab2.reset_counte_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_4_LC_11_11_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_4_LC_11_11_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.shifter_4_LC_11_11_4 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \buart.Z_rx.shifter_4_LC_11_11_4  (
            .in0(_gnd_net_),
            .in1(N__6506),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6181),
            .ce(N__6072),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.de0.g0_5_LC_11_11_5 .C_ON=1'b0;
    defparam \Glue_Lab2.de0.g0_5_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.de0.g0_5_LC_11_11_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Glue_Lab2.de0.g0_5_LC_11_11_5  (
            .in0(_gnd_net_),
            .in1(N__5119),
            .in2(_gnd_net_),
            .in3(N__5488),
            .lcout(),
            .ltout(\Glue_Lab2.de0.g0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.de0.g0_9_LC_11_11_6 .C_ON=1'b0;
    defparam \Glue_Lab2.de0.g0_9_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.de0.g0_9_LC_11_11_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Glue_Lab2.de0.g0_9_LC_11_11_6  (
            .in0(N__5455),
            .in1(N__5176),
            .in2(N__5392),
            .in3(N__5384),
            .lcout(),
            .ltout(\Glue_Lab2.g0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.reset_count_RNO_0_3_LC_11_11_7 .C_ON=1'b0;
    defparam \Glue_Lab2.reset_count_RNO_0_3_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.reset_count_RNO_0_3_LC_11_11_7 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \Glue_Lab2.reset_count_RNO_0_3_LC_11_11_7  (
            .in0(N__5304),
            .in1(N__6685),
            .in2(N__5260),
            .in3(N__5257),
            .lcout(\Glue_Lab2.reset_counte_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_2_LC_11_12_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_2_LC_11_12_0 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.shifter_2_LC_11_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_2_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6613),
            .lcout(bu_rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6187),
            .ce(N__6071),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_5_LC_11_12_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_5_LC_11_12_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.shifter_5_LC_11_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_5_LC_11_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5131),
            .lcout(bu_rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6187),
            .ce(N__6071),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_fast_4_LC_11_12_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_4_LC_11_12_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.shifter_fast_4_LC_11_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_fast_4_LC_11_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6519),
            .lcout(buart__rx_shifter_fast_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6187),
            .ce(N__6071),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_tx_data_RNO_1_5_LC_11_13_0 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_tx_data_RNO_1_5_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.Gl_tx_data_RNO_1_5_LC_11_13_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Glue_Lab2.Gl_tx_data_RNO_1_5_LC_11_13_0  (
            .in0(_gnd_net_),
            .in1(N__6031),
            .in2(_gnd_net_),
            .in3(N__6007),
            .lcout(),
            .ltout(\Glue_Lab2.g0_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.Gl_tx_data_RNO_0_5_LC_11_13_1 .C_ON=1'b0;
    defparam \Glue_Lab2.Gl_tx_data_RNO_0_5_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.Gl_tx_data_RNO_0_5_LC_11_13_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Glue_Lab2.Gl_tx_data_RNO_0_5_LC_11_13_1  (
            .in0(N__5983),
            .in1(N__5953),
            .in2(N__5923),
            .in3(N__5920),
            .lcout(\Glue_Lab2.Gl_subtract_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.S_0_s_ac0_5_0_0_LC_11_13_3 .C_ON=1'b0;
    defparam \Lab_UT.S_0_s_ac0_5_0_0_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.S_0_s_ac0_5_0_0_LC_11_13_3 .LUT_INIT=16'b1111100010000000;
    LogicCell40 \Lab_UT.S_0_s_ac0_5_0_0_LC_11_13_3  (
            .in0(N__5883),
            .in1(N__5814),
            .in2(N__5662),
            .in3(N__5733),
            .lcout(\Lab_UT.S_0_s_ac0_5_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.S_1_c3_c_LC_11_13_5 .C_ON=1'b0;
    defparam \Lab_UT.S_1_c3_c_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.S_1_c3_c_LC_11_13_5 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \Lab_UT.S_1_c3_c_LC_11_13_5  (
            .in0(N__5884),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5815),
            .lcout(),
            .ltout(\Lab_UT.S_1_c3_cZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.S_1_c4_LC_11_13_6 .C_ON=1'b0;
    defparam \Lab_UT.S_1_c4_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.S_1_c4_LC_11_13_6 .LUT_INIT=16'b1000000011101010;
    LogicCell40 \Lab_UT.S_1_c4_LC_11_13_6  (
            .in0(N__5734),
            .in1(N__5677),
            .in2(N__5665),
            .in3(N__5660),
            .lcout(),
            .ltout(\Lab_UT.C_out41_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.L2_led_1_4_LC_11_13_7 .C_ON=1'b0;
    defparam \Lab_UT.L2_led_1_4_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.L2_led_1_4_LC_11_13_7 .LUT_INIT=16'b0000111111101110;
    LogicCell40 \Lab_UT.L2_led_1_4_LC_11_13_7  (
            .in0(N__5593),
            .in1(N__5587),
            .in2(N__5575),
            .in3(N__5572),
            .lcout(led_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_12_8_0 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_12_8_0 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_12_8_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_2_LC_12_8_0  (
            .in0(_gnd_net_),
            .in1(N__6877),
            .in2(_gnd_net_),
            .in3(N__6909),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6184),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_12_8_1 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_12_8_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_12_8_1 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_3_LC_12_8_1  (
            .in0(N__6910),
            .in1(N__6821),
            .in2(N__6885),
            .in3(N__6857),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6184),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_8_LC_12_10_1 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_8_LC_12_10_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.shifter_8_LC_12_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \buart.Z_tx.shifter_8_LC_12_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6764),
            .lcout(\buart.Z_tx.shifterZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6183),
            .ce(N__6701),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.de0.g0_8_LC_12_11_1 .C_ON=1'b0;
    defparam \Glue_Lab2.de0.g0_8_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.de0.g0_8_LC_12_11_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Glue_Lab2.de0.g0_8_LC_12_11_1  (
            .in0(N__6675),
            .in1(N__6596),
            .in2(N__6529),
            .in3(N__6472),
            .lcout(\Glue_Lab2.g0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.sDelay.delayReg_3_LC_12_12_0 .C_ON=1'b0;
    defparam \Lab_UT.sDelay.delayReg_3_LC_12_12_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.sDelay.delayReg_3_LC_12_12_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Lab_UT.sDelay.delayReg_3_LC_12_12_0  (
            .in0(N__6307),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6373),
            .lcout(\Lab_UT.sDelay.delayRegZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6191),
            .ce(),
            .sr(_gnd_net_));
    defparam \Glue_Lab2.de0.g0_6_LC_12_12_5 .C_ON=1'b0;
    defparam \Glue_Lab2.de0.g0_6_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \Glue_Lab2.de0.g0_6_LC_12_12_5 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Glue_Lab2.de0.g0_6_LC_12_12_5  (
            .in0(N__6679),
            .in1(N__6612),
            .in2(N__6528),
            .in3(N__6473),
            .lcout(\Glue_Lab2.g0_8_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.sDelay.delayReg_2_LC_12_12_6 .C_ON=1'b0;
    defparam \Lab_UT.sDelay.delayReg_2_LC_12_12_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.sDelay.delayReg_2_LC_12_12_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Lab_UT.sDelay.delayReg_2_LC_12_12_6  (
            .in0(N__6306),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6382),
            .lcout(\Lab_UT.sDelay.delayRegZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6191),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.sDelay.delayReg_4_LC_12_12_7 .C_ON=1'b0;
    defparam \Lab_UT.sDelay.delayReg_4_LC_12_12_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.sDelay.delayReg_4_LC_12_12_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.sDelay.delayReg_4_LC_12_12_7  (
            .in0(_gnd_net_),
            .in1(N__6367),
            .in2(_gnd_net_),
            .in3(N__6308),
            .lcout(L2_adder_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6191),
            .ce(),
            .sr(_gnd_net_));
endmodule // latticehx1k
